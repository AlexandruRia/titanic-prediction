���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.0�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJ�
hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h4�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh(�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M�nodes�h*h-K ��h/��R�(KM��h4�V64�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h}hLK ��h~hLK��hhLK��h�h]K��h�h]K ��h�hLK(��h�h]K0��h�h4�u1�����R�(Kh8NNNJ����J����K t�bK8��uK@KKt�b�B@E         �                     @"��p�?�           8�@               u                    �?.y0��k�?�            �s@ u r n        "                    �?Hث3���?�            @m@ 497e131                           �?     ��?)             P@5.3"}1                         0�FF@�'N��?&            �N@ hHbQ                           s�,@�q�����?             9@        ������������������������       �                     @�5bQ         	                 �܅3@8�A�0��?             6@ iHbQ  ������������������������       �                     @        
                        p�i@@�\��N��?             3@                                  �?��
ц��?	             *@                                   �?      �?             @        ������������������������       �                     �?                                  �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �<@և���X�?             @ }4bQ  ������������������������       �                     @Pq4bQ  ������������������������       �                     @�g4bQ                             �?�q�q�?             @s4bQ  ������������������������       �                     @�t4bQ  ������������������������       �                      @�x4bQ                             �?�����H�?             B@z4bQ  ������������������������       �                     9@�{4bQ                          p"�X@���|���?             &@}4bQ                            �8@؇���X�?             @ s4bQ  ������������������������       �                     �? O4bQ  ������������������������       �                     @ [4bQ                             �?      �?             @ b4bQ  ������������������������       �                     �?�GbQ  ������������������������       �                     @ GbQ          !                    �?�q�q�?             @GbQ  ������������������������       �                      @��aQ  ������������������������       �                     �?��aQ  #       &                   �9@���Q��?i            @e@        $       %                    �?��s����?             5@        ������������������������       �                     @i
aQ  ������������������������       �                     1@.�aQ  '       f                  x#J@p�B<F]�?[            �b@�aQ  (       G                     �?��c`��?L            �^@      0@)       >                   �>@8����?              G@�aQ  *       +                    �?��
ц��?             :@ �aQ  ������������������������       �                     @      @,       -                   �<@�q�q�?             5@ aQ  ������������������������       �                     @      �?.       =                    R@�<ݚ�?             2@�aQ  /       0                 03:@@�0�!��?             1@      @������������������������       �                     @��aQ  1       <                   �J@���!pc�?	             &@�aQ  2       3                 03k:@      �?              @ �aQ  ������������������������       �                     �?      @4       ;                    H@����X�?             @�aQ  5       :                 X��B@r�q��?             @     �?6       7                 `fF<@      �?             @ �aQ  ������������������������       �                      @9�aQ  8       9                 �|Y=@      �?              @ �aQ  ������������������������       �                     �?<�aQ  ������������������������       �                     �?��aQ  ������������������������       �                      @��aQ  ������������������������       �                     �?      @������������������������       �                     @       @������������������������       �                     �?'�aQ  ?       @                 `f~I@ףp=
�?             4@�aQ  ������������������������       �                     (@G�aQ  A       B                 `��I@      �?              @      �?������������������������       �                     �?6aQ  C       D                 03�I@؇���X�?             @ �aQ  ������������������������       �                     �?b�aQ  E       F                    �?r�q��?             @      �?������������������������       �                     �?PaQ  ������������������������       �                     @       @H       e                    >@&:~�Q�?,             S@"aQ  I       X                    �?�Y�R_�?+            �Q@ "aQ  J       K                   @B@ �o_��?             9@ (aQ  ������������������������       �                     "@��aQ  L       S                    -@     ��?             0@�aQ  M       P                   �'@      �?              @ -aQ  N       O                   �J@      �?              @ �aQ  ������������������������       �                     �?faQ  ������������������������       �                     �?       Q       R                    D@�q�q�?             @ aQ  ������������������������       �                     @��aQ  ������������������������       �                      @NaQ  T       W                   �H@      �?              @�aQ  U       V                   �E@      �?             @ haQ  ������������������������       �                      @�LaQ  ������������������������       �                      @��aQ  ������������������������       �                     @!^aQ  Y       d                    �?���}<S�?             G@aQ  Z       c                   @A@��-�=��?            �C@ �aQ  [       b                   �@@������?
             1@aQ  \       ]                 �|Y=@�r����?	             .@ aQ  ������������������������       �                     @:�aQ  ^       _                   �'@�<ݚ�?             "@aQ  ������������������������       �                     @8BaQ  `       a                 �|�=@�q�q�?             @ �aQ  ������������������������       �                      @        ������������������������       �                     �?NaQ  ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     @��aQ  ������������������������       �                     @f�aQ  g       t                 03�U@PN��T'�?             ;@�aQ  h       i                    <@��s����?             5@ �aQ  ������������������������       �                     @^KaQ  j       k                    ?@      �?	             0@        ������������������������       �                     �??�aQ  l       m                    B@z�G�z�?             .@ =aQ  ������������������������       �                     @�aaQ  n       o                    C@�z�G��?             $@ aQ  ������������������������       �                      @�%aQ  p       q                    �?      �?              @ &aQ  ������������������������       �                     @�aQ  r       s                 0� Q@      �?             @ �aQ  ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    :@���B���?3            �S@ �aQ  ������������������������       �        
             1@9�aQ  x                          �8@�jTM��?)            �N@ �aQ  y       ~                    @�g�y��?             ?@ �aQ  z       {                 ��W@      �?             @        ������������������������       �                      @�aQ  |       }                 �(\�?      �?              @ aQ  ������������������������       �                     �?5)aQ  ������������������������       �                     �?��aQ  ������������������������       �                     ;@H9aQ  �       �                    �?��S���?             >@�aQ  �       �                  DT@�ՙ/�?             5@       �       �                     �?�n_Y�K�?	             *@        �       �                 X�,D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       �       �                 �UA@r�q��?             @       �       �                   @A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�~�@
�?�            �x@        �       �                    7@�g�y��?             ?@        �       �                 03�@ףp=
�?             $@       ������������������������       �                     "@       ������������������������       �                     �?        ������������������������       �                     5@        �       
                ��Y7@�?��+�?�             w@       �       �                    /@����I�?�            �t@        �       �                    $@      �?             8@       ������������������������       �        	             .@       �       �                 �&�)@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       �       �                    �?����Y��?�            s@        �       �                    �?���ȫ�?/            �T@        �       �                    �?�MI8d�?            �B@       �       �                    �?      �?             @@       ������������������������       �                     6@       �       �                  S�-@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @       �       �                 `�@1@z�G�z�?             @       ������������������������       �                     @       ������������������������       �                     �?        �       �                     @X�<ݚ�?            �F@       �       �                  s@~�4_�g�?             F@        ������������������������       �                     @        �       �                   �3@      �?             D@        ������������������������       �                     �?        �       �                   �4@�99lMt�?            �C@        ������������������������       �                     @        �       �                 ��/@b�2�tk�?             B@       �       �                    �?�z�G��?             >@       �       �                   �5@�û��|�?             7@        ������������������������       �                     �?        �       �                    �?���|���?             6@       �       �                   P&@�q�q�?             5@       �       �                 �|�;@�z�G��?             4@       �       �                 pf�@�n_Y�K�?             *@        ������������������������       �                      @        �       �                 pf� @���!pc�?             &@       �       �                   �9@և���X�?             @       �       �                   �6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��� @؇���X�?             @       ������������������������       �                     @        �       �                  SE"@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@�@+��?�            �k@        �       �                    �?�<ݚ�?             2@       �       �                   @@$�q-�?
             *@        �       �                 �|�:@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     "@        �       �                   �2@���Q��?             @        ������������������������       �                      @       ������������������������       �                     @       �       �                    �?�M��?}            �i@        �       �                    �?XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        �       �                 �?�@h�V���?l             f@        �       �                   �?@�k~X��?.             R@       ������������������������       �        %             L@        �       �                   @@@      �?	             0@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     ,@        �       �                   �1@�ջ����?>             Z@        ������������������������       �                     (@        �       	                   �?��H�?7             W@       �                          �?z�G�z�?2            @U@       �       �                 @3�@*�s���?1             U@        �       �                   �?@      �?             ,@        �       �                   �9@�q�q�?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �A@      �?              @        ������������������������       ��q�q�?             @       ������������������������       ����Q��?             @        �       �                   �2@؇���X�?*            �Q@        ������������������������       �                     @        �       �                 ��) @pH����?)            �P@        �       �                   �3@ 7���B�?             ;@        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   �9@R���Q�?             D@        ������������������������       �                     1@        �                          (@��+7��?             7@       �                          ?@���Q��?             .@                              �|Y=@      �?              @        ������������������������       �                     @                              �̜!@���Q��?             @        ������������������������       �                     �?                              �|�=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                              ��T?@��-�=��?            �C@       ������������������������       �                     9@                                 �?����X�?             ,@        ������������������������       �                     @                                 @���|���?             &@                                @���Q��?             $@                             ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�b�values�h*h-K ��h/��R�(KMKK��h]�BP        {@     Pq@     �`@      f@      ^@     �\@      2@      G@      1@      F@      *@      (@              @      *@      "@      @              $@      "@      @      @      @      @      �?               @      @              @       @              @      @              @      @              @       @      @                       @      @      @@              9@      @      @      �?      @      �?                      @      @      �?              �?      @              �?       @               @      �?             �Y@      Q@      1@      @              @      1@             @U@      P@     @T@     �D@      @@      ,@      ,@      (@              @      ,@      @              @      ,@      @      ,@      @      @               @      @      @      @              �?      @       @      @      �?      @      �?       @              �?      �?      �?                      �?       @                      �?      @                      �?      2@       @      (@              @       @              �?      @      �?      �?              @      �?              �?      @             �H@      ;@     �H@      6@      @      2@              "@      @      "@      @      @      �?      �?              �?      �?              @       @      @                       @       @      @       @       @               @       @                      @      E@      @     �A@      @      *@      @      *@       @      @              @       @      @              �?       @               @      �?                       @      6@              @                      @      @      7@      @      1@              @      @      (@      �?              @      (@              @      @      @       @              �?      @              @      �?      @              @      �?                      @      .@     �O@              1@      .@      G@      �?      >@      �?      @               @      �?      �?              �?      �?                      ;@      ,@      0@       @      *@       @      @      @      �?              �?      @              @      @              @      @                       @      @      @      �?       @      �?                       @      @      �?      @      �?              �?      @               @             �r@      Y@      >@      �?      "@      �?      "@                      �?      5@             �p@     �X@     @m@     �W@      @      5@              .@      @      @              @      @      �?       @              �?      �?      �?                      �?     �l@     �R@      ?@     �I@      @      ?@       @      >@              6@       @       @       @                       @      @      �?      @                      �?      9@      4@      9@      3@              @      9@      .@              �?      9@      ,@      @              6@      ,@      5@      "@      ,@      "@              �?      ,@       @      ,@      @      ,@      @       @      @               @       @      @      @      @      @      �?              �?      @                       @      @              @      �?      @              �?      �?              �?      �?                      �?              �?      @              �?      @      �?                      @              �?      i@      7@      ,@      @      (@      �?      @      �?       @              �?      �?      "@               @      @       @                      @     @g@      3@      <@      �?      <@                      �?     �c@      2@     �Q@      �?      L@              .@      �?      �?      �?              �?      �?              ,@             �U@      1@      (@             �R@      1@      Q@      1@     �P@      1@      @      @       @      @       @       @       @                       @               @      @      @       @      �?      @       @      N@      $@              @      N@      @      :@      �?              �?      :@              A@      @      1@              1@      @      "@      @       @      @              @       @      @              �?       @       @       @                       @      @               @              �?              @             �A@      @      9@              $@      @      @              @      @      @      @       @      @              @       @              @              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ/��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @���*1�?�           8�@                                   @�7����?            �G@     "@                            �?Pa�	�?            �@@      @                           �?z�G�z�?             @        ������������������������       �                     �?       @������������������������       �                     @      9@������������������������       �                     <@      @       	                 ��T?@؇���X�?             ,@       @������������������������       �                      @        
                           @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               z                     @��?a�?�           ��@               !                    �?V$�݆��?�            �r@                                 0Cd=@Pns��ޭ?O            �`@                                  @E@$Q�q�?"            �O@                               ���*@p���?             I@ �� ���                        `f�)@�IєX�?	             1@ f4bQ  ������������������������       �                     (@ m4bQ                             :@z�G�z�?             @ /aQ                             5@      �?              @ �aQ  ������������������������       �                     �?�s4bQ  ������������������������       �                     �?�u4bQ  ������������������������       �                     @ w4bQ  ������������������������       �                    �@@��aQ                             �?�θ�?             *@:aQ                          ���;@ףp=
�?             $@{4bQ  ������������������������       �                     "@UHaQ  ������������������������       �                     �?�~4bQ                             �?�q�q�?             @  GbQ  ������������������������       �                      @�GbQ  ������������������������       �                     �?laQ  ������������������������       �        -            �Q@GbQ  "       y                    �?4>���?t             e@�FbQ  #       8                 `ff:@�{��?��?n            @d@ �aQ  $       '                    5@ >�֕�?0            �Q@ aQ  %       &                   �2@      �?              @ aQ  ������������������������       �                     �?��FbQ  ������������������������       �                     �?�aQ  (       )                 �|Y=@ =[y��?.             Q@ �aQ  ������������������������       �                     4@T�aQ  *       7                   �*@      �?#             H@�aQ  +       ,                 `f�)@ȵHPS!�?             :@�aQ  ������������������������       �                     0@;�aQ  -       .                 �|�=@�z�G��?             $@      @������������������������       �                     �?��aQ  /       4                   @D@�<ݚ�?             "@�aQ  0       3                   �A@؇���X�?             @ �aQ  1       2                    @@�q�q�?             @ �FbQ  ������������������������       �                      @T�aQ  ������������������������       �                     �?      <@������������������������       �                     @��aQ  5       6                   �G@      �?              @ �aQ  ������������������������       �                     �?��aQ  ������������������������       �                     �?�aQ  ������������������������       �                     6@K�aQ  9       V                    �?�)
;&��?>             W@ �aQ  :       U                     �?�e����?            �C@�aQ  ;       T                   �H@��J�fj�?            �B@�aQ  <       Q                   @C@�g�y��?             ?@�aQ  =       >                   �4@�û��|�?             7@ �aQ  ������������������������       �                     @5�aQ  ?       P                 �̾w@�G�z��?             4@�FbQ  @       M                    �?ҳ�wY;�?             1@�aQ  A       D                 �|�;@�q�q�?
             (@ �aQ  B       C                 Ȉ�P@�q�q�?             @
      ������������������������       �                      @respondi������������������������       �                     �?�4aQ  E       L                   �A@�<ݚ�?             "@\aQ  F       K                 ��2>@�q�q�?             @ r   rG       H                 `f&;@�q�q�?             @  aQ  ������������������������       �                     �?�}t|I       J                 ���<@      �?              @ "aQ  ������������������������       �                     �?OaQ  ������������������������       �                     �? aQ  ������������������������       �                     @4FaQ  ������������������������       �                     @ bound_hN       O                   �7@���Q��?             @ YaQ  ������������������������       �                      @ ound af������������������������       �                     @��aQ  ������������������������       �                     @�aQ  R       S                 ���X@      �?              @+aQ  ������������������������       �                     @    ����������������������������       �                     �?naQ  ������������������������       �                     @ �aQ  ������������������������       �                      @�0aQ  W       f                  i?@�c�����?"            �J@ 
X       e                   @>@p�ݯ��?             3@>aQ  Y       d                   �J@�t����?
             1@}}nZ       c                 `f�;@X�<ݚ�?             "@}n|[       ^                 �|�?@����X�?             @ |t�\       ]                 �|�<@      �?              @ aQ  ������������������������       �                     �?}&d||#������������������������       �                     �?  us�|_       `                   �C@z�G�z�?             @ �aQ  ������������������������       �                     @KaQ  a       b                    H@      �?              @ }.}/d������������������������       �                     �?}5|�d������������������������       �                     �?  }6t������������������������       �                      @|8��������������������������       �                      @|: }"������������������������       �                      @{�aQ  g       x                     �?@�0�!��?             A@|<< |h       i                   �A@�n`���?             ?@ �aQ  ������������������������       �                     "@*haQ  j       w                    �?���!pc�?             6@�aQ  k       v                    �?����X�?             5@�aQ  l       m                   �B@�z�G��?             4@ �aQ  ������������������������       �                     @b0aQ  n       u                 `f�K@@�0�!��?             1@r6   r7o       p                   �C@��S�ۿ?             .@$aQ  ������������������������       �                     "@ �aQ  q       r                    �?r�q��?             @ naQ  ������������������������       �                     @JrI   Zs       t                  x#J@      �?              @ undr  ������������������������       �                     �?_reduct������������������������       �                     �?.aQ  ������������������������       �                      @ step_fr������������������������       �                     �?��aQ  ������������������������       �                     �?�aQ  ������������������������       �                     @M�aQ  ������������������������       �                     @5aQ  {       �                   �@@\�Yf�?�            �v@�aQ  |       �                    �?�8a�ME�?�            �s@ �aQ  }       �                    �?@��Pl3�?<            @X@ �aQ  ~       �                    �?     ��?             @@vaQ         �                    �?�>4և��?             <@  rX   �       �                    �?�IєX�?             1@ �aQ  ������������������������       �                      @        �       �                 �|�6@��S�ۿ?
             .@  aQ  ������������������������       �                     @0aQ  �       �                 ���@�8��8��?             (@ �aQ  ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?���|���?             &@        �       �                   �,@z�G�z�?             @        ������������������������       �                     �? aQ  ������������������������       �                     @�aQ  ������������������������       �                     @        ������������������������       �                     @�aQ  �       �                    �?&����?(            @P@       �       �                 03�-@>���Rp�?%             M@       �       �                    �?�LQ�1	�?             G@       �       �                    �?8�Z$���?             :@       �       �                 ���@r�q��?             8@ ,aQ  ������������������������       �                     "@        �       �                   @@������?             .@       �       �                   �5@�q�q�?             "@        ������������������������       �                     �?�aQ  �       �                 �|=@      �?              @ vaQ  ������������������������       �                      @       �       �                 �|�=@�q�q�?             @ aQ  ������������������������       �      �?             @        ������������������������       �                      @�aQ  �       �                 �|Y=@r�q��?             @        ������������������������       �                     �? |aQ  ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y;@ףp=
�?             4@ kaQ  ������������������������       �                     �?       �       �                  s�@�KM�]�?             3@        ������������������������       �                     @ �aQ  �       �                    �?؇���X�?
             ,@       ������������������������       �8�Z$���?	             *@        ������������������������       �                     �?       �       �                 ��.@�q�q�?             (@ �aQ  ������������������������       �                     @        �       �                 ��$1@և���X�?             @        ������������������������       �                     @        �       �                   �2@      �?             @ ?aQ  ������������������������       �                     �?       ������������������������       �                     @�aQ  ������������������������       �                     @        �       �                    �?�nYU}�?�             k@	aQ  �       �                    @�C�F��?o            �e@FaQ  �       �                 �|�=@�R����?n            �e@       �       �                    �?*~k���?b            �b@        �       �                  s@�eP*L��?             6@ �aQ  ������������������������       �                     @?aQ  �       �                    4@�q�q�?             2@ �aQ  �       �                    �?      �?             @        ������������������������       �                     @'aQ  ������������������������       �                     �?        �       �                 �|�;@d}h���?
             ,@saQ  �       �                 pff@ףp=
�?             $@        �       �                   �7@      �?              @ �aQ  ������������������������       �                     �? �aQ  ������������������������       �                     �?        ������������������������       �                      @	aQ  �       �                    �?      �?             @aQ  ������������������������       �                      @�aQ  ������������������������       �                      @ �aQ  �       �                    �?x�]AgȽ?T             `@       �       �                    �?`Jj��?R             _@       �       �                 ���@�IєX�?N            �]@ �aQ  �       �                   �5@����X�?             @ �aQ  ������������������������       �                     @       �       �                 �&b@      �?             @       ������������������������       �                      @ �aQ  ������������������������       �                      @ DaQ  �       �                   �0@���>4ֵ?I             \@ aQ  �       �                 pFD!@      �?             @        ������������������������       �      �?              @ �aQ  ������������������������       �                      @        �       �                 @3�!@ 7���B�?E             [@3aQ  �       �                 @3�@������?6            �T@�aQ  �       �                 �?$@���J��?!            �I@ 7aQ  �       �                 ��@���N8�?             5@       ������������������������       �        	             1@        �       �                 �|Y8@      �?             @        ������������������������       �                     �?       ������������������������       ��q�q�?             @ �aQ  ������������������������       �                     >@ saQ  �       �                 pf� @��a�n`�?             ?@EaQ  �       �                   �4@�8��8��?             8@ �aQ  �       �                   �2@����X�?             @        ������������������������       �                      @2aQ  �       �                 0S5 @���Q��?             @�aQ  ������������������������       ��q�q�?             @�aQ  ������������������������       �                      @ �aQ  ������������������������       �                     1@ �aQ  �       �                    8@؇���X�?             @iaQ  ������������������������       �                     @        ������������������������       �                     �?��aQ  ������������������������       �                     :@       �       �                 �Y�@z�G�z�?             @ eaQ  ������������������������       �                      @       �       �                 pF�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @ 4aQ  ������������������������       �                     @       �       �                   @@@8�A�0��?             6@�aQ  �       �                    �?      �?
             2@       �       �                    �?     ��?	             0@        ������������������������       �                     @        �       �                   �?@��
ц��?             *@ 6aQ  ������������������������       �                     @       �       �                 d�6@@���Q��?             $@       �       �                 ��I @և���X�?             @aQ  �       �                 P�@      �?             @ eaQ  ������������������������       �                      @       ������������������������       �      �?              @       ������������������������       �                     @�aQ  ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @ �aQ  ������������������������       �                      @       �       �                 �̜2@d}h���?             E@ aQ  �       �                    <@�	j*D�?             *@�aQ  �       �                 P�@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@paQ  ������������������������       �                      @       ������������������������       �                     =@�aQ  ������������������������       �                     H@        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �{@     �p@      *@      A@      �?      @@      �?      @      �?                      @              <@      (@       @       @              @       @      @                       @     �z@     �m@     �a@     @d@      @      `@      @     �M@      �?     �H@      �?      0@              (@      �?      @      �?      �?              �?      �?                      @             �@@      @      $@      �?      "@              "@      �?               @      �?       @                      �?             �Q@      a@     �@@      `@     �@@     �P@      @      �?      �?      �?                      �?     @P@      @      4@             �F@      @      7@      @      0@              @      @              �?      @       @      @      �?       @      �?       @                      �?      @              �?      �?              �?      �?              6@             �O@      =@      7@      0@      5@      0@      .@      0@      ,@      "@      @              &@      "@      &@      @       @      @      �?       @               @      �?              @       @      @       @      �?       @              �?      �?      �?      �?                      �?      @              @              @       @               @      @                      @      �?      @              @      �?              @               @              D@      *@      (@      @      (@      @      @      @       @      @      �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?       @               @                       @      <@      @      9@      @      "@              0@      @      .@      @      ,@      @              @      ,@      @      ,@      �?      "@              @      �?      @              �?      �?      �?                      �?               @      �?              �?              @              @             �q@     �R@     �m@     �R@      N@     �B@      "@      7@      @      7@      �?      0@               @      �?      ,@              @      �?      &@      �?                      &@      @      @      @      �?              �?      @                      @      @             �I@      ,@      F@      ,@      D@      @      6@      @      4@      @      "@              &@      @      @      @              �?      @       @       @              @       @       @       @       @              @      �?              �?      @               @              2@       @      �?              1@       @      @              (@       @      &@       @      �?              @       @              @      @      @      @              �?      @      �?                      @      @             `f@      C@     @b@      =@     @b@      ;@     �`@      2@      (@      $@              @      (@      @      �?      @              @      �?              &@      @      "@      �?      �?      �?              �?      �?               @               @       @       @                       @     @^@       @      ]@       @      \@      @      @       @      @               @       @       @                       @     �Z@      @      @      �?      �?      �?       @              Z@      @     �S@      @      I@      �?      4@      �?      1@              @      �?      �?               @      �?      >@              <@      @      6@       @      @       @       @              @       @      �?       @       @              1@              @      �?      @                      �?      :@              @      �?       @               @      �?              �?       @              @              *@      "@      "@      "@      @      "@              @      @      @      @              @      @      @      @      �?      @               @      �?      �?      @                      @       @              @                       @     �@@      "@      @      "@       @      "@       @                      "@       @              =@              H@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJu�7hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�F         D                    �?���Yb�?�           8�@    -
         )                    �?&ջ�{��?]            @b@9/bQ                             �?JJ����?;            �W@      @                           �?��hJ,�?             A@    @j@������������������������       �                     ;@       @                        �ܙH@����X�?             @     9@������������������������       �                     @      @������������������������       �                      @       @	       
                   �2@      �?'             N@        ������������������������       �                     @                                     @����>4�?$             L@                                  @B@�ՙ/�?             5@                               ���<@      �?             0@        ������������������������       �                     @                                   �?�n_Y�K�?	             *@                               03SA@���Q��?             $@        ������������������������       �                     @                                @�6M@և���X�?             @      ;@������������������������       �                     @      "@                        X�,@@      �?             @                               �|Y<@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?       @������������������������       �                      @       @                        �nc@�q�q�?             @        ������������������������       �                     �?      1@                        �̾w@      �?              @      (@������������������������       �                     �?      @������������������������       �                     �?        ������������������������       �                     @      G@       "                 �|Y=@�#-���?            �A@      �?        !                   @@z�G�z�?             $@     0@������������������������       �                      @      (@������������������������       �                      @      @#       $                 ���@`2U0*��?             9@ �EbQ  ������������������������       �                     &@�HbQ  %       (                 �|�=@@4և���?
             ,@HbQ  &       '                   @@      �?              @     0@������������������������       �r�q��?             @p�EbQ  ������������������������       �                      @�5bQ  ������������������������       �                     @p�EbQ  *       3                     @R�}e�.�?"             J@�EbQ  +       ,                    �?z�G�z�?             >@�EbQ  ������������������������       �                     4@0�EbQ  -       2                    �?���Q��?             $@     �?.       1                     �?�q�q�?             @�EbQ  /       0                 �U�X@z�G�z�?             @�EbQ  ������������������������       �                     @��EbQ  ������������������������       �                     �?      @������������������������       �                     �?0�EbQ  ������������������������       �                     @       4       =                    �?���|���?
             6@ �EbQ  5       <                    �?և���X�?             ,@�GbQ  6       9                    �?�eP*L��?             &@ �EbQ  7       8                   �-@և���X�?             @ �EbQ  ������������������������       �                     @��EbQ  ������������������������       �                     @p�EbQ  :       ;                 �|Y3@      �?             @ �GbQ  ������������������������       �                     @��EbQ  ������������������������       �                     �?05bQ  ������������������������       �                     @��EbQ  >       C                 03�-@      �?              @�EbQ  ?       B                    �?�q�q�?             @      @@       A                 �&�)@      �?              @ �EbQ  ������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @      @E                       `f�S@��f
a�?r           ��@       F       �                 `f�$@�K�7���?]           Ȁ@        G       \                    �?��1��?�            �n@        H       S                   �6@�g�y��?             ?@        I       R                    �?r�q��?
             (@       J       O                    �?�<ݚ�?             "@       K       L                    �?؇���X�?             @        ������������������������       �                      @        M       N                   �3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       Q                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       Y                 ��@�d�����?             3@        U       V                 ���@�q�q�?             @        ������������������������       �                     �?        W       X                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       [                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ]       b                   �0@d��]a��?�            �j@        ^       _                 pf�@���!pc�?             &@        ������������������������       �                     @        `       a                 pFD!@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        c       l                    �?����p�?�            �i@        d       e                 ���@�>4և��?             <@        ������������������������       �                      @        f       g                 �|Y=@      �?
             4@        ������������������������       �                     @        h       k                 X��A@�t����?	             1@       i       j                    �?؇���X�?             ,@       ������������������������       �8�Z$���?             *@        ������������������������       �                     �?        ������������������������       �                     @        m       �                 �|�=@����!p�?u             f@       n       {                 �?$@ ,V�ނ�?V            �_@        o       x                 ���@�L���?            �B@       p       q                     @�g�y��?             ?@        ������������������������       �                     "@        r       s                  Md@���7�?             6@        ������������������������       �                     &@        t       u                    7@�C��2(�?             &@        ������������������������       �                     @        v       w                   �8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                 �|�;@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        |       �                    �?�x�E~�?;            @V@       }       �                    �?`���i��?:             V@       ~                        @3�@�D�e���?8            @U@        ������������������������       �                    �C@        �       �                   �;@�nkK�?             G@       �       �                   �9@�>����?             ;@910,15.�       �                   �3@ ��WV�?             :@ 58,,S
6�       �                   �2@�C��2(�?             &@ 0.5,,S
������������������������       �                     @ rgue)",�       �                 0S5 @؇���X�?             @ iss. El������������������������       �      �?              @,"Ander������������������������       �                     @ale,39,������������������������       �        	             .@,,0,0,S������������������������       �                     �?  Jane",������������������������       �                     3@e,,0,0,������������������������       �                     @ male,35������������������������       �                     �? 24,1,2,�       �                   @@@ףp=
�?             I@ 1,1,347�       �                 �?�@�	j*D�?             *@ K Stanl������������������������       �                     @ss. Mar�       �                    ?@X�<ݚ�?             "@ r. Lawr�       �                 �̌!@      �?              @ oni",ma������������������������       �                     �? son Jr"������������������������       �                     �?id",male�       �                 ��I @և���X�?             @ard",ma������������������������       ����Q��?             @  ""Dai"������������������������       �                      @ick",mal�       �                      @�?�|�?            �B@ les Leo������������������������       �                     @. Gretch�       �                   �C@г�wY;�?             A@ndyeff,�       �                   @C@�IєX�?             1@nnell, ������������������������       �        
             .@orth, Mr������������������������       �      �?              @,3,"Lun������������������������       �        	             1@ 3,1,1,"�       �                    �?��c���?�            0r@ 34,0,1,�       �                    �?ڷv���?I            �\@ ,0,3,"S�       �                    �?Hm_!'1�?            �H@ avis, M������������������������       �                     �? Mr. Ant�       �                    �?      �?             H@,"Colly�       �                     @ �Cc}�?             <@Panula,�       �                     �?$�q-�?             :@ .6875,,������������������������       �                     @6.1,,S
�       �                   �A@�C��2(�?             6@2,,S
64�       �                   �9@�IєX�?
             1@ B35,C
6�       �                   �'@؇���X�?             @ 8,27.9,������������������������       �                     @ 5,1,3,"�       �                   �3@      �?              @ 46,1,1,������������������������       �                     �? D33,C
6������������������������       �                     �? 48,1,1,������������������������       �                     $@35.5,A26�       �                   �D@z�G�z�?             @ .55,,S
������������������������       �                     �? A. 2314������������������������       �                     @958,,S
�       �                 ��&@      �?              @ 653,0,3������������������������       �                     �?,,S
654������������������������       �                     �?,7.8292������������������������       �                     4@0,36522�       �                     @8�A�0��?*            �P@ ,S.O.C.�       �                     �?�}�+r��?             3@ 349223,������������������������       �                     @32,1,1,�       �                    �?��S�ۿ?             .@ e,23,0,�       �                    B@      �?             @8,0,2,3������������������������       �                     @ ",male,������������������������       �                     �?e,40,0,������������������������       �        	             &@ ,47,0,0�       �                    �?��k=.��?            �G@ 0,34921������������������������       �                      @,1,0,ST�       �                   @1@���V��?            �F@ e,32,2,�       �                    �?���|���?             &@on",mal�       �                    D@����X�?             @",male,�       �                 �|�;@      �?             @ 0,A/5 3������������������������       �                      @ummins W������������������������       �                      @ Thomas ������������������������       �                     @ ,29750,�       �                    0@      �?             @ 2750,52������������������������       �                      @ C.A. 24������������������������       �                      @244270,1�       �                    @l��\��?             A@ 6,0,,S
�       �                    @����X�?             @12,7.77������������������������       �                     @ 0,34282������������������������       �                      @0,4138,9�       �                    @ 7���B�?             ;@",femal������������������������       �                     7@ ke Mart�       �                   @D@      �?             @ ,"Peter������������������������       �                     �?ssab, Mr������������������������       �                     @ vigen, �                          �?��|���?t             f@dwin, M�       �                    �?H%u��?T            @_@ rown, M�       �                    �?      �?              @2,"Laro������������������������       �                     @ 2123,41������������������������       �                     �?3101295,�       �                 `fF:@�S#א��?N            @]@,10.170�       �                    4@����p�?+             Q@ 0,35003�       �                    &@�<ݚ�?             "@ emale,1������������������������       �                      @ n",male������������������������       �                     @e,4,0,1�       �                     @����˵�?$            �M@56.4958�       �                   �*@���.�6�?             G@695,0,1�       �                 `f�)@ܷ��?��?             =@ hapman,������������������������       �                     @Kelly, M�       �                   �A@�LQ�1	�?             7@ss. Kat�       �                    @@d}h���?             ,@ayer, M������������������������       �                      @,"Humbl������������������������       �      �?             @ .65,F G������������������������       �                     "@ Force)"������������������������       �                     1@thorne,������������������������       �                     *@ 03,0,3,�                         �Q@Jm_!'1�?#            �H@,0,3,"G�                          �?r�q��?"             H@,"Hanse�                             @t/*�?!            �G@"Morley�       �                   �;@"pc�
�?             F@ 50655,2�       �                    �?�q�q�?             @ 0,0,223������������������������       �                     �?male,42,�       �                    7@      �?              @ ,female������������������������       �                     �?  Gonios������������������������       �                     �?,"Mayne,�       �                   �>@�p ��?            �D@ ,0,PC 1�       �                    K@     ��?             0@,113028�       �                   `G@�eP*L��?             &@1,0,199�       �                   @>@      �?              @,0,0,75�       �                 `f�;@؇���X�?             @250647,�       �                 �|�<@      �?             @ ",male,������������������������       �                     �?e Louis������������������������       �                     @ Miss. E������������������������       �                     @ 19,0,3,������������������������       �                     �?ohnson, ������������������������       �                     @,"Harper������������������������       �                     @722,0,3�       �                  x#J@`2U0*��?             9@
723,0,������������������������       �                     1@724,0,2�       �                 `�iJ@      �?              @ ,1,"Cha������������������������       �                     �? 726,0,3������������������������       �                     @ ,2,"Ren������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��[�8��?             �I@                                +@J�8���?             =@        ������������������������       �                     $@        ������������������������       �                     3@                                 @���7�?             6@       	      
                   �?      �?
             0@       ������������������������       �                     *@                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�>4և��?             <@                                M@H%u��?             9@                              �k@�8��8��?             8@                               @E@�nkK�?             7@       ������������������������       �                     3@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �}@     �m@      P@     �T@      I@      F@      @      =@              ;@      @       @      @                       @     �F@      .@              @     �F@      &@      *@       @       @       @      @              @       @      @      @              @      @      @      @              �?      @      �?      �?              �?      �?                       @      �?       @              �?      �?      �?      �?                      �?      @              @@      @       @       @       @                       @      8@      �?      &@              *@      �?      @      �?      @      �?       @              @              ,@      C@      @      8@              4@      @      @       @      @      �?      @              @      �?              �?              @               @      ,@      @       @      @      @      @      @      @                      @      @      �?      @                      �?              @       @      @       @      �?      �?      �?              �?      �?              �?                      @     �y@     @c@     `y@     ``@     �j@     �@@      0@      .@       @      $@       @      @      �?      @               @      �?      @      �?                      @      �?      �?              �?      �?                      @      ,@      @       @      @      �?              �?      @              @      �?              (@      �?              �?      (@             �h@      2@       @      @      @              @      @              @      @             �g@      .@      7@      @       @              .@      @              @      .@       @      (@       @      &@       @      �?              @             �d@      $@     @^@      @      A@      @      >@      �?      "@              5@      �?      &@              $@      �?      @              @      �?              �?      @              @       @      @              �?       @     �U@       @     �U@       @     �T@       @     �C@              F@       @      9@       @      9@      �?      $@      �?      @              @      �?      �?      �?      @              .@                      �?      3@              @              �?             �F@      @      "@      @      @              @      @      �?      �?      �?                      �?      @      @       @      @       @              B@      �?      @             �@@      �?      0@      �?      .@              �?      �?      1@              h@     �X@     �E@      R@      @     �F@      �?              @     �F@      @      9@       @      8@              @       @      4@      �?      0@      �?      @              @      �?      �?      �?                      �?              $@      �?      @      �?                      @      �?      �?      �?                      �?              4@     �C@      ;@      �?      2@              @      �?      ,@      �?      @              @      �?                      &@      C@      "@               @      C@      @      @      @      @       @       @       @       @                       @      @               @       @               @       @              ?@      @      @       @      @                       @      :@      �?      7@              @      �?              �?      @             �b@      :@     �[@      .@      @      �?      @                      �?     �Y@      ,@     �O@      @      @       @               @      @              L@      @     �E@      @      :@      @      @              4@      @      &@      @       @              @      @      "@              1@              *@              D@      "@      D@       @     �C@       @      B@       @      �?       @              �?      �?      �?      �?                      �?     �A@      @      &@      @      @      @      @       @      @      �?      @      �?              �?      @              @                      �?              @      @              8@      �?      1@              @      �?              �?      @              @              �?                      �?      D@      &@      3@      $@              $@      3@              5@      �?      .@      �?      *@               @      �?       @                      �?      @              @      7@      @      6@       @      6@      �?      6@              3@      �?      @              @      �?              �?              �?               @      �?       @                      �?�t�bub�$>     hhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��!XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         l                 ��%@�*���?�           8�@      =@                           /@,PY��?�             v@  u r n ������������������������       �                     @      @                        ���@j�q����?�            �u@ �aQ  ������������������������       �                    �E@��aQ         3                 P�*@�A��t��?�            0s@ �aQ         2                 �|Y>@J��D��?A             [@"5bQ         1                    �?���Q �?8            �X@�aQ  	       
                 ��@r�qG�?7             X@ f2bQ  ������������������������       �                     �?���XQ                             �?�|R���?6            �W@ a4bQ                            �3@���B���?             :@ ��XQ                          �?@�q�q�?             @ ��[Q  ������������������������       �                     �?�r�aQ  ������������������������       �                      @���XQ                             �?�LQ�1	�?             7@��XQ                             8@�C��2(�?             6@      @������������������������       �                     "@      .@                        ��@8�Z$���?	             *@      @                        ���@�C��2(�?             &@      �?                           �?�q�q�?             @      @������������������������       �                      @      @������������������������       �                     �?        ������������������������       �                      @      @                           @      �?              @      @������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                     �?      �?       $                   �<@�㙢�c�?&            @Q@      �?       #                   �6@�C��2(�?            �@@                                  �3@�S����?
             3@       @������������������������       �                      @       @!       "                    �?���!pc�?             &@      &@������������������������       �                     @      �?������������������������       �                      @        ������������������������       �                     ,@      @%       .                    �?      �?             B@     @&       '                 ���@z�G�z�?             9@       @������������������������       �                      @      �?(       )                 �|Y=@�t����?             1@        ������������������������       �                     �?       @*       +                 ���@      �?
             0@      @������������������������       ����Q��?             @      @,       -                 �Y�@�C��2(�?             &@      ;@������������������������       �                     @      @������������������������       �      �?              @      @/       0                 ��,@���|���?             &@       ������������������������       �                     @       @������������������������       ��q�q�?             @       @������������������������       �                      @       @������������������������       �        	             $@        4       i                    �?ȭ^���?x            �h@     �?5       <                 �?�@��ɉ�?v            `h@      �?6       ;                 �̌@�L#���?)            �P@       @7       8                 �|Y=@���y4F�?             3@       ������������������������       �        
             *@      �?9       :                 ��]@�q�q�?             @      �?������������������������       �                      @      "@������������������������       �                     @      @������������������������       �                     H@      @=       B                     @     ��?M             `@      @>       A                   �J@�+e�X�?             9@     "@?       @                    �?�����?             3@      "@������������������������       �                     @        ������������������������       �                     *@      �?������������������������       �                     @6aQ  C       N                 @3�@�v�G���??            �Y@ �aQ  D       G                    �?      �?             0@ �aQ  E       F                   �9@���Q��?             @     �?������������������������       �                     @PaQ  ������������������������       �                      @       @H       I                    :@���|���?             &@ "aQ  ������������������������       �                     @ "aQ  J       K                   �?@և���X�?             @ (aQ  ������������������������       �                     �?��aQ  L       M                   �A@      �?             @ �aQ  ������������������������       �      �?              @ -aQ  ������������������������       �      �?             @ �aQ  O       V                   �:@�=C|F�?4            �U@ aQ  P       U                   �3@`Ӹ����?            �F@        Q       T                 0S5 @�����?
             5@ aQ  R       S                   �1@�q�q�?             @ �aQ  ������������������������       �                     �?NaQ  ������������������������       �                      @�aQ  ������������������������       �                     2@ haQ  ������������������������       �                     8@�LaQ  W       X                   �;@d}h���?             E@ �aQ  ������������������������       �                     @!^aQ  Y       h                   �?@8�Z$���?            �C@aQ  Z       [                 ��) @      �?             8@�aQ  ������������������������       �        	             &@aQ  \       ]                   �<@��
ц��?             *@ aQ  ������������������������       �                     @:�aQ  ^       c                 P�*"@���Q��?             $@ aQ  _       `                 pf� @z�G�z�?             @ BaQ  ������������������������       �                      @ �aQ  a       b                    �?�q�q�?             @        ������������������������       �                      @NaQ  ������������������������       �                     �?        d       e                 ���"@���Q��?             @        ������������������������       �                      @��aQ  f       g                 �|Y=@�q�q�?             @ �aQ  ������������������������       �                      @�aQ  ������������������������       �                     �? �aQ  ������������������������       �        	             .@^KaQ  j       k                   �#@      �?             @        ������������������������       �                      @?�aQ  ������������������������       �                      @ =aQ  m       �                  x#J@��d���?�            Pv@aaQ  n       �                    �?~���n��?�            Pp@ aQ  o       �                    @t�I��n�?R            @]@%aQ  p       u                    @f�����?N            �[@ &aQ  q       r                    @�}�+r��?             3@�aQ  ������������������������       �        
             0@ �aQ  s       t                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       �                     @ �&�T�?B             W@�aQ  w       �                   �H@�j��b�?(            �M@�aQ  x       �                    �?,�+�C�?%            �K@�aQ  y       z                     �?<���D�?            �@@ �aQ  ������������������������       �                     @        {       �                   �7@8�Z$���?             :@�aQ  |       �                    �?������?             .@aQ  }       �                    :@d}h���?             ,@ )aQ  ~                           �?      �?             @ �aQ  ������������������������       �                      @H9aQ  ������������������������       �                      @�aQ  �       �                    �?ףp=
�?	             $@        ������������������������       �                     �?        �       �                   �*@�����H�?             "@       �       �                 `f�)@؇���X�?             @        ������������������������       �                     �?        �       �                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     6@        �       �                 03�9@      �?             @       ������������������������       �                      @       ������������������������       �                      @        �       �                    �?4���C�?            �@@       �       �                 ��.@\X��t�?             7@       �       �                    �?�	j*D�?
             *@        �       �                 �|Y6@և���X�?             @       �       �                   �,@      �?             @        ������������������������       �                      @       �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @       �       �                   �*@r�q��?             @        ������������������������       �                     �?       ������������������������       �                     @       �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 �|Y>@r�q��?             @        ������������������������       �                     @        �       �                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       �       �                 ���0@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@       ������������������������       �                     @       �       �                    @�q�q�?g             b@       �       �                    !@�θ�?^            @`@        ������������������������       �                     $@        �       �                 �&@r�q��?W             ^@        ������������������������       �                     �?       �       �                     �?�?��,�?V            �]@        �       �                 ��";@���j��?             G@        �       �                 ��$:@և���X�?
             ,@        ������������������������       �                     @        �       �                   �J@���!pc�?             &@       �       �                   @G@�����H�?             "@       �       �                    D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @       ������������������������       �                      @       �       �                    �?     ��?             @@       �       �                 ���=@�����?             5@        ������������������������       �                     $@       �       �                 p�i@@"pc�
�?             &@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                  �>@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @        �       �                   �<@���!pc�?	             &@        ������������������������       �                      @        �       �                 �|Y>@�����H�?             "@        �       �                 �|Y=@      �?             @        ������������������������       �                     �?       �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                     @        �       �                   �*@�F��O�?8            @R@        �       �                   �@@�㙢�c�?             7@       ������������������������       �        
             (@        �       �                   �)@���|���?	             &@        ������������������������       �                      @        �       �                   �A@X�<ݚ�?             "@        ������������������������       �      �?             @        �       �                   @D@z�G�z�?             @        ������������������������       �                      @       �       �                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`2U0*��?%             I@       �       �                 ��.@`Ql�R�?"            �G@        �       �                     @$�q-�?
             *@        ������������������������       �                     @       �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        �                          @     ��?B             X@       �       �                    �?�n`���??            @W@       �       �                   �5@f>�cQ�?-            �N@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @       �       �                    �?$�q-�?'             J@       �       �                      @�IєX�?&            �I@       �       �                   �B@ �q�q�?#             H@       �       �                    �?�IєX�?             A@       ������������������������       �                     <@        �       �                    �?�q�q�?             @       �       �                 X�,@@      �?             @       �       �                 p"�b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     �?                                �7@     ��?             @@                                 �?�C��2(�?             &@                                �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�ՙ/�?             5@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       `|@     p@     �q@     �P@              @     �q@     �O@     �E@             �n@     �O@     �R@      A@      P@      A@      O@      A@              �?      O@     �@@      @      5@       @      �?              �?       @              @      4@       @      4@              "@       @      &@      �?      $@      �?       @               @      �?                       @      �?      �?      �?                      �?      �?             �L@      (@      >@      @      0@      @       @               @      @              @       @              ,@              ;@      "@      4@      @       @              (@      @              �?      (@      @       @      @      $@      �?      @              @      �?      @      @      @               @      @       @              $@             @e@      =@      e@      ;@     �O@      @      .@      @      *@               @      @       @                      @      H@             @Z@      7@      3@      @      *@      @              @      *@              @             �U@      1@      $@      @      @       @      @                       @      @      @      @              @      @              �?      @      @      �?      �?       @       @      S@      &@     �E@       @      3@       @      �?       @      �?                       @      2@              8@             �@@      "@              @     �@@      @      2@      @      &@              @      @      @              @      @      �?      @               @      �?       @               @      �?              @       @       @              �?       @               @      �?              .@               @       @               @       @             �d@     �g@     @b@     �\@      @@     @U@      :@     @U@      �?      2@              0@      �?       @      �?                       @      9@     �P@      @     �J@      @     �I@      @      =@              @      @      6@      @      &@      @      &@       @       @               @       @              �?      "@              �?      �?       @      �?      @              �?      �?      @              @      �?                       @      �?                      &@              6@       @       @               @       @              3@      ,@      $@      *@      "@      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?              �?      @              �?      "@              @      �?      @              @      �?      �?      �?                      �?      "@      �?              �?      "@              @             �\@      >@      Y@      >@              $@      Y@      4@              �?      Y@      3@     �@@      *@      @       @      @              @       @      �?       @      �?      @               @      �?       @              @       @              ;@      @      3@       @      $@              "@       @      �?       @              �?      �?      �?      �?                      �?       @               @      @               @       @      �?      @      �?      �?               @      �?              �?       @              @             �P@      @      3@      @      (@              @      @       @              @      @      �?      @      @      �?       @               @      �?              �?       @              H@       @      G@      �?      (@      �?      @              @      �?      @              �?      �?      �?                      �?      A@               @      �?              �?       @              ,@              5@     �R@      2@     �R@      "@      J@      @      @              @      @              @      H@      @      H@       @      G@       @      @@              <@       @      @      �?      @      �?      �?              �?      �?                       @      �?      �?              �?      �?                      ,@      �?       @              �?      �?      �?      �?                      �?      �?              "@      7@      �?      $@      �?      @      �?                      @              @       @      *@              *@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJC�NhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         p                     @���%&�?�           8�@ d4bQ         '                 �|Y=@N�ec�?�            ps@      @       
                 ��*@"��$�?G            �[@      5@       	                    �?      �?             8@      4@                           �?"pc�
�?             &@�aQ                          `f�)@�<ݚ�?             "@�aQ  ������������������������       �                     @"5bQ  ������������������������       �                      @�aQ  ������������������������       �                      @        ������������������������       �        
             *@               "                 `fmj@�N��D�?6            �U@                                  �?���(\��?2             T@                                  6@�C��2(�?)            �P@                                   9@���|���?             &@       ������������������������       �                     @                                   �?z�G�z�?             @        ������������������������       �                     �?      @������������������������       �                     @      .@                           �?h㱪��?#            �K@      @������������������������       �                    �B@      �?                            �?�����H�?
             2@     @                           5@��S�ۿ?             .@      @������������������������       �                     �?        ������������������������       �                     ,@      @                           �?�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @                                   �?d}h���?	             ,@     �?                            �?�����H�?             "@      �?������������������������       �                     �?       ������������������������       �                      @       @        !                    �?���Q��?             @      @������������������������       �                     @      &@������������������������       �                      @      �?#       &                 0U�o@և���X�?             @       $       %                    5@z�G�z�?             @      @������������������������       �                     �?     @������������������������       �                     @       @������������������������       �                      @      �?(       9                    �?4��@���?�             i@        )       ,                    �?�nkK�?1            @Q@       @*       +                 03�=@`2U0*��?             9@      @������������������������       �                     �?      @������������������������       �                     8@      ;@-       6                    L@���7�?             F@     @.       /                   �B@��Y��]�?            �D@     @������������������������       �                     8@       0       5                    -@�IєX�?             1@       @1       2                   �'@�q�q�?             @       @������������������������       �                     �?       @3       4                    D@      �?              @        ������������������������       �                     �?     �?������������������������       �                     �?      �?������������������������       �        	             ,@       @7       8                   �L@�q�q�?             @        ������������������������       �                     �?      �?������������������������       �                      @      �?:       o                   �J@��ׂ�?Z            ``@     "@;       n                 p�w@������?F            @Z@     @<       a                   �G@��z6��?D             Y@     @=       >                   �)@� ���?6            @S@      @������������������������       �        	             ,@     "@?       `                   �F@��s����?-            �O@     "@@       [                    �?�T`�[k�?(            �J@       A       L                    �?��Q���?             D@      @B       K                    �?     ��?
             0@       C       J                    C@�q�q�?	             .@       D       I                 ��2>@����X�?             ,@        E       H                 ���<@      �?              @       F       G                 ��";@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        M       Z                    �?      �?             8@       N       W                   @D@���!pc�?             6@       O       V                 `f�<@@�0�!��?             1@       P       U                 `fF:@���!pc�?             &@       Q       T                 `fv3@z�G�z�?             $@       R       S                 �|�=@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                     �?���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                      @        \       ]                   �B@$�q-�?             *@        ������������������������       �                     @        ^       _                 03�U@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        b       c                 `f4@
;&����?             7@        ������������������������       �                     @        d       i                    �?     ��?	             0@        e       f                    �?�q�q�?             @        ������������������������       �                      @        g       h                 ���X@      �?             @       ������������������������       �                      @        ������������������������       �                      @        j       k                 ���E@ףp=
�?             $@       ������������������������       �                      @        l       m                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        q                          @z6�>��?            y@       r       s                 ���@�o6�
�?�            �x@        ������������������������       �                     ;@        t                          @.�6�G,�?�             w@       u       �                    �?H?�߽��?�            �v@        v       �                    �?�\��N��?H            �\@        w       |                    �?,���i�?            �D@       x       {                 ���@      �?             @@        y       z                 0��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        }       ~                    @X�<ݚ�?             "@        ������������������������       �                      @               �                  S�2@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                      @       �       �                 ���&@�q�q�?             @ (aQ  ������������������������       �                     �?�8aQ  �       �                 �|Y=@      �?              @ �aQ  ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @       �       �                    @:PZ(8?�?-            @R@        �       �                    @z�G�z�?             @ aQ  ������������������������       �                      @��aQ  �       �                    @�q�q�?             @        ������������������������       �                     �?��aQ  ������������������������       �                      @       �       �                    ,@�t����?)             Q@        ������������������������       �                     $@        �       �                   �"@J�8���?$             M@        �       �                    @�ՙ/�?             5@4aQ  �       �                    ;@���Q��?             4@       �       �                    �?������?
             .@       �       �                 pf� @d}h���?	             ,@       �       �                   �7@�C��2(�?             &@ �aQ  ������������������������       �                     @�}aQ  �       �                 �&B@z�G�z�?             @        ������������������������       �                     �?�aQ  ������������������������       �                     @       �       �                    3@�q�q�?             @ �aQ  ������������������������       �                     �?        ������������������������       �                      @��aQ  ������������������������       �                     �?        �       �                 �?� @z�G�z�?             @       ������������������������       �                     @}saQ  ������������������������       �                     �?       ������������������������       �                     �?        �       �                 03�1@��G���?            �B@�aQ  �       �                    �?�X����?             6@       �       �                     @ҳ�wY;�?             1@       �       �                   �3@������?
             .@        ������������������������       �                     �?�aQ  �       �                   �0@d}h���?	             ,@       �       �                 �|�;@8�Z$���?             *@        ������������������������       �                      @        �       �                 ���.@���Q��?             @GaQ  �       �                    �?      �?             @       �       �                   �@@      �?              @ �aQ  ������������������������       �                     �?       ������������������������       �                     �?0aQ  ������������������������       �                      @�MaQ  ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @^�aQ  �       �                   �;@z�G�z�?             @ GaQ  ������������������������       �                     �?ɪaQ  ������������������������       �                     @        ������������������������       �                     .@�.aQ  �       �                 ��@H%u��?�            @o@        ������������������������       �                     @f{aQ  �       �                    #@0�v����?�            �n@        �       �                     @     ��?             0@ �aQ  ������������������������       �                     @��aQ  �       �                    @ףp=
�?             $@       �       �                    �?z�G�z�?             @ aQ  ������������������������       �                     �?�#aQ  �       �                 ���A@      �?             @ �aQ  �       �                    @      �?              @ �aQ  ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @�aQ  ������������������������       �                     @b�aQ  �       �                    �?,���>�?�            �l@        �       �                 03�-@д>��C�?'             M@       �       �                 �|Y=@ףp=
�?              I@ �aQ  �       �                   �<@�<ݚ�?             "@KaQ  ������������������������       �                     @"aQ  ������������������������       �                      @        �       �                 �|Y?@��p\�?            �D@�aQ  �       �                    �?ܷ��?��?             =@       �       �                 ���@�����H�?             ;@ ;aQ  ������������������������       �                     @�aQ  �       �                 P�J@؇���X�?             5@>aQ  �       �                 ���@R���Q�?             4@        �       �                    �?�����H�?             "@       ������������������������       �r�q��?             @       ������������������������       �                     @       ������������������������       �"pc�
�?             &@H�aQ  ������������������������       �                     �?7{aQ  ������������������������       �                      @�LaQ  ������������������������       �                     (@��aQ  �       �                 ��.@      �?              @        ������������������������       �                     @�aQ  �       �                    �?���Q��?             @ �aQ  ������������������������       �                     �?2�aQ  �       �                    �?      �?             @�aQ  ������������������������       �                     @8�aQ  ������������������������       �                     �?�paQ  �                         @@@���y�?p            �e@       �                          �?D��*�4�?\            @a@�aQ  �                          �?�[|x��?U            �_@       �       �                 �!&B@�H�@=��?M            �[@maQ  �       �                 �|�=@ �h�7W�?J            �Z@       �       �                 @3�@��8�$>�?C            @X@       ������������������������       �        $             H@       �       �                 @�!@Hm_!'1�?            �H@;aQ  �       �                   � @PN��T'�?             ;@       �       �                 0S5 @�r����?             .@�aQ  �       �                   �3@؇���X�?             ,@        �       �                    1@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @�=aQ  ������������������������       �                     &@        ������������������������       �                     �?       �       �                   �7@r�q��?             (@%aQ  ������������������������       �                      @�laQ  �       �                 �|Y<@      �?             @        ������������������������       �                      @        ������������������������       �                      @t�aQ  ������������������������       �                     6@       �       �                   �?@�<ݚ�?             "@       �       �                   �>@���Q��?             @ �aQ  �       �                 �̌!@      �?              @        ������������������������       �                     �?SaQ  ������������������������       �                     �?<�aQ  �       �                 pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?oxaQ  ������������������������       �                     @        �       �                    ;@z�G�z�?             @ �aQ  ������������������������       �                      @                                  >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     (@        ������������������������       �                    �A@                               �:@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       �{@     �p@     �`@      f@      <@     �T@      .@      "@       @      "@       @      @              @       @                       @      *@              *@     �R@      "@     �Q@      @      N@      @      @              @      @      �?              �?      @               @     �J@             �B@       @      0@      �?      ,@      �?                      ,@      �?       @      �?                       @      @      &@      �?       @      �?                       @       @      @              @       @              @      @      @      �?              �?      @                       @     �Z@     �W@      @     �P@      �?      8@      �?                      8@       @      E@      �?      D@              8@      �?      0@      �?       @              �?      �?      �?      �?                      �?              ,@      �?       @      �?                       @     �Y@      <@     @S@      <@     @S@      7@     @P@      (@      ,@             �I@      (@     �D@      (@      =@      &@      &@      @      $@      @      $@      @      @      @      @      �?              �?      @                      @      @                      �?      �?              2@      @      0@      @      ,@      @       @      @       @       @      @       @               @      @              @                      �?      @               @      @      �?      �?      �?       @       @              (@      �?      @              @      �?      @                      �?      $@              (@      &@      @              @      &@      @       @       @               @       @               @       @              �?      "@               @      �?      �?      �?                      �?              @      :@             0s@     @W@     �r@     @W@      ;@             0q@     @W@      q@     �V@      K@      N@      @      B@      �?      ?@      �?       @               @      �?                      =@      @      @               @      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                       @     �H@      8@      �?      @               @      �?       @      �?                       @      H@      4@      $@              C@      4@       @      *@       @      (@      @      &@      @      &@      �?      $@              @      �?      @      �?                      @       @      �?              �?       @              �?              @      �?      @                      �?              �?      >@      @      .@      @      &@      @      &@      @              �?      &@      @      &@       @       @              @       @      @      �?      �?      �?              �?      �?               @                      �?              �?               @      @      �?              �?      @              .@             �k@      >@              @     �k@      ;@      "@      @              @      "@      �?      @      �?      �?              @      �?      �?      �?      �?                      �?       @              @             `j@      4@      H@      $@     �F@      @      @       @      @                       @      C@      @      :@      @      8@      @      @              2@      @      1@      @       @      �?      @      �?      @              "@       @      �?               @              (@              @      @              @      @       @              �?      @      �?      @                      �?     `d@      $@      `@      $@      ]@      $@     @Y@      $@      Y@      @     @W@      @      H@             �F@      @      7@      @      *@       @      (@       @      �?       @      �?                       @      &@              �?              $@       @       @               @       @               @       @              6@              @       @      @       @      �?      �?      �?                      �?       @      �?       @                      �?      @              �?      @               @      �?       @      �?                       @      .@              (@             �A@              �?      @              @      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�R�[hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         \                    �?�s�ˈ.�?�           8�@    -
         U                 p�H@�d�����?�            �l@              4                    �?Ҙ$�Ų�?k            �d@     @                            @�<ݚ�?=            �X@ �aQ         
                    �?�(\����?             D@

    N                          �J@�nkK�?             7@       ������������������������       �                     4@ �a]Q         	                 `f�2@�q�q�?             @ where u������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@                                   �?:���W�?#            �M@                                   �?�+e�X�?             9@                                H�%@���Q��?             $@        ������������������������       �                     @                                03�-@z�G�z�?             @        ������������������������       �                     @      @                        �|Y=@      �?              @      .@������������������������       �                     �?      @������������������������       �                     �?      �?                        X�,A@�r����?             .@     @������������������������       �                     *@      @������������������������       �                      @               /                    �?�ʻ����?             A@     @       .                    �?*;L]n�?             >@     @                           '@П[;U��?             =@       @������������������������       �                     @                                  �4@      �?             :@      �?������������������������       �                     @      �?       )                 `��!@\X��t�?             7@              (                    C@������?	             .@      @        !                 P�@d}h���?             ,@       @������������������������       �                     @      �?"       '                 �|Y>@      �?              @     8@#       &                 �|�;@      �?             @       $       %                   �8@      �?              @      4@������������������������       �                     �?      &@������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @      �?������������������������       �                     �?      @*       +                    ;@      �?              @      @������������������������       �                     @      �?,       -                   �@@�q�q�?             @      �?������������������������       �                      @      �?������������������������       �                     �?      @������������������������       �                     �?      �?0       1                    @      �?             @      �?������������������������       �                     �?        2       3                 ��l4@�q�q�?             @       @������������������������       �                     �?      @������������������������       �                      @      @5       <                     @�'�=z��?.            �P@       @6       9                    6@؇���X�?             5@      @7       8                 ��m1@      �?             @      �?������������������������       �                      @      $@������������������������       �                      @      @:       ;                   �B@�IєX�?             1@      @������������������������       �                     0@       @������������������������       �                     �?        =       @                    �?f.i��n�?            �F@        >       ?                 ��.@�q�q�?             @        ������������������������       �                      @      �?������������������������       �                     @       @A       J                 03�1@��Sݭg�?            �C@        B       I                    �?�q�q�?             (@       C       H                 ��Y.@���Q��?             $@       D       G                    �?z�G�z�?             @       E       F                    6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        K       P                    @�>����?             ;@       L       O                 ���4@���7�?             6@        M       N                 03C3@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             3@        Q       R                 ��T?@z�G�z�?             @        ������������������������       �                      @        S       T                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        V       [                 ���Q@$Q�q�?+            �O@        W       X                    �?�J�4�?             9@       ������������������������       �                     3@        Y       Z                 ���P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     C@        ]       �                    �?���A�
�?*           0~@        ^       k                 ��K.@N��c��?1            @S@        _       d                   �6@������?            �D@        `       a                    �?      �?             @        ������������������������       �                     �?        b       c                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                 �|=@�?�|�?            �B@        ������������������������       �                     &@        g       j                   @@ ��WV�?             :@       h       i                 ���@�C��2(�?             &@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     .@        l       w                    �?b�2�tk�?             B@       m       r                 �|Y<@�z�G��?             4@        n       q                    9@����X�?             @        o       p                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        s       v                   �F@$�q-�?
             *@        t       u                 X�,@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        x                           �?      �?             0@       y       |                 ��G@և���X�?
             ,@        z       {                 ��3@      �?              @        ������������������������       �                     @        ������������������������       �                     @        }       ~                 ���X@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �/@|g�&��?�            `y@, Mr. N�       �                    �?<N_�U��?�            �p@�GbQ  �       �                 �?�@     �?�             p@ �GbQ  �       �                     @������?M            �^@ GbQ  ������������������������       �                     &@ McMahon�       �                    �?�h����?E             \@ r. Frid�       �                  ��@8�Z$���?             *@ Miss. A������������������������       �                      @ r. Joha�       �                    �?"pc�
�?	             &@9GbQ  �       �                 �|Y=@�<ݚ�?             "@ GbQ  ������������������������       �                     �?ns, Mrs.�       �                 ��(@      �?              @GbQ  ������������������������       �r�q��?             @ )",fema������������������������       �                      @ayden",������������������������       �                      @ ,male,2�       �                   �7@��:x�ٳ?:            �X@ en Mony������������������������       �                     A@��GbQ  �       �                 �Yu@����?&            @P@n, Mr. �       �                 �&B@(N:!���?            �A@. Victo�       �                   �8@`Jj��?             ?@ Joseph �       �                 �&b@���Q��?             @ �FbQ  ������������������������       �                     @��GbQ  ������������������������       �                      @O2. 310������������������������       �                     :@�$GbQ  �       �                    �?      �?             @ 31945,1������������������������       �                      @ GbQ  ������������������������       �                      @ nnerstr������������������������       �                     >@�aGbQ  �       �                   �0@���H��?N            �`@ 2,"Navr�       �                 �̌!@�q�q�?             @ 080,26,������������������������       �                      @��GbQ  ������������������������       �                     �? 0,S.O.P�       �                   �*@ ����?L            @`@e)",fem�       �                   �A@���5��?D            �\@�FbQ  �       �                   �<@8�Z$���?7            �V@ Blyler�       �                   �3@$�q-�?             J@ Martin"�       �                     @������?	             .@ rles Du�       �                    &@      �?             @ <8bQ  ������������������������       �      �?              @"Corn, M������������������������       �                      @ iljanic�       �                   �1@���!pc�?             &@ ter. Th������������������������       �                     @0�GbQ  �       �                 0S5 @և���X�?             @  James ������������������������       �                     @�FbQ  ������������������������       �                     @47068,7������������������������       �                    �B@ .GbQ  �       �                 ��)"@��Sݭg�?            �C@�GbQ  �       �                   �?@�KM�]�?             3@kie""",�       �                   �>@8�Z$���?             *@h Marth�       �                 �|Y=@�8��8��?
             (@ �FbQ  ������������������������       �                     �?��GbQ  �       �                 ��) @�C��2(�?	             &@�0bQ  ������������������������       �                     "@an der �       �                 pf� @      �?              @ �GbQ  ������������������������       �                     �?son, Mi������������������������       �                     �?��GbQ  ������������������������       �                     �? ,,S
175������������������������       �                     @58bQ  �       �                 �|�=@���Q��?             4@ ?8bQ  ������������������������       �                     @7,,S
17�       �                   �@@�t����?             1@-GbQ  �       �                    $@�θ�?	             *@ =GbQ  �       �                   �?@      �?             @ �FbQ  ������������������������       �                     @`�FbQ  ������������������������       �                     �? 3,"Aspl������������������������       �                     "@ 875,,S
������������������������       �      �?             @@�6bQ  ������������������������       �                     7@��FbQ  ������������������������       �                     0@ 7,50,A3�       �                    �?���|���?             &@frey)",�       �                     @X�<ݚ�?             "@ 5bQ  ������������������������       �                     �?0�GbQ  �       �                   �*@      �?              @ <GbQ  �       �                 xFT$@���Q��?             @ Rosa)",������������������������       �                      @0
GbQ  ������������������������       �                     @ Christi������������������������       �                     @�GbQ  ������������������������       �                      @`GbQ  �       �                    @4kMU*m�?X            `a@ �GbQ  �       �                   �;@������?             .@ 146.520������������������������       �                     @.75,,Q
1�       �                    @      �?              @ 9,8.404������������������������       �                     @,0,0,37������������������������       �                     @0GbQ  �                          �?���b��?P             _@5bQ  �       �                    �? �&�T�?:             W@5bQ  �       �                     @���3�E�?$             J@88bQ  �       �                 ��$:@�*/�8V�?             �G@ ,male,4������������������������       �        	             .@�8GbQ  �       �                   �>@      �?             @@�FbQ  �       �                 `fF<@�t����?             1@�FbQ  �       �                    K@      �?             $@GbQ  �       �                 03k:@����X�?             @ [3bQ  ������������������������       �                     �?�\GbQ  �       �                 �|�<@�q�q�?             @ ,24,0,0������������������������       �                      @��FbQ  �       �                 X��B@      �?             @ hn Henr������������������������       �                     �?`�GbQ  �       �                   @G@�q�q�?             @lip",ma������������������������       �      �?              @female,������������������������       �                     �?a",fema������������������������       �                     @@�GbQ  ������������������������       �                     @ s. Albi������������������������       �                     .@0 GbQ  �       �                 �|�>@���Q��?             @ Victor�       �                 �T�C@�q�q�?             @ acken, ������������������������       �                     �? George�       �                 �|�;@      �?              @ �GbQ  ������������������������       �                     �?Maxfiel������������������������       �                     �? Ivar S������������������������       �                      @0IGbQ  �       �                    �?      �?             D@[GbQ  �       �                  x#J@r٣����?            �@@ahlstro������������������������       �        
             1@bre, Mi�       �                    F@      �?             0@�GbQ  �       �                 `f�K@�q�q�?             (@75,C83,�       �                    7@      �?              @ .775,,S������������������������       �                     @`GbQ  �       �                 `�iJ@z�G�z�?             @ 077,31.������������������������       �                      @�,GbQ  �       �                    @@�q�q�?             @ �FbQ  ������������������������       �                      @ ,44,1,0������������������������       �                     �?,female������������������������       �                     @ �GbQ  ������������������������       �                     @ Henry",�       �                 �|�:@����X�?             @ �FbQ  ������������������������       �                     @erine ""                            @�q�q�?             @ . Regin������������������������       �                     �?        ������������������������       �                      @                                 @      �?             @@                                �?`Jj��?             ?@                                 @�X�<ݺ?             2@        ������������������������       �                     @              
                   @@4և���?	             ,@             	                   0@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �|@     @o@      N@      e@      L@     @[@      6@     @S@      �?     �C@      �?      6@              4@      �?       @      �?                       @              1@      5@      C@      @      3@      @      @              @      @      �?      @              �?      �?              �?      �?               @      *@              *@       @              .@      3@      *@      1@      *@      0@              @      *@      *@      @              $@      *@      @      &@      @      &@              @      @      @      @      �?      �?      �?      �?                      �?       @                      @      �?              @       @      @              �?       @               @      �?                      �?       @       @              �?       @      �?              �?       @              A@      @@      @      2@       @       @               @       @              �?      0@              0@      �?              ?@      ,@       @      @       @                      @      =@      $@      @       @      @      @      @      �?      @      �?              �?      @              �?                      @               @      9@       @      5@      �?       @      �?       @                      �?      3@              @      �?       @               @      �?              �?       @              @     �M@      @      5@              3@      @       @               @      @                      C@     y@     �T@     �M@      2@     �B@      @      �?      @              �?      �?       @               @      �?              B@      �?      &@              9@      �?      $@      �?      @              @      �?      .@              6@      ,@      ,@      @       @      @       @      �?       @                      �?              @      (@      �?      @      �?      @                      �?       @               @       @      @       @      @      @              @      @              �?      @              @      �?               @             `u@      P@      n@      :@     @m@      6@     @]@      @      &@             �Z@      @      &@       @       @              "@       @      @       @              �?      @      �?      @      �?       @               @             �W@      @      A@             �N@      @      ?@      @      =@       @      @       @      @                       @      :@               @       @               @       @              >@             @]@      0@      �?       @               @      �?              ]@      ,@      Y@      ,@     @S@      ,@      H@      @      &@      @      @      �?      �?      �?       @               @      @      @              @      @              @      @             �B@              =@      $@      1@       @      &@       @      &@      �?      �?              $@      �?      "@              �?      �?              �?      �?                      �?      @              (@       @              @      (@      @      $@      @      �?      @              @      �?              "@               @       @      7@              0@              @      @      @      @              �?      @      @       @      @       @                      @      @               @             @Y@      C@      @      &@              @      @      @              @      @             @X@      ;@     �P@      9@     �B@      .@     �A@      (@      .@              4@      (@      @      (@      @      @       @      @              �?       @      @               @       @       @      �?              �?       @      �?      �?              �?      @                      @      .@               @      @       @      �?      �?              �?      �?              �?      �?                       @      >@      $@      9@       @      1@               @       @      @       @      @      @      @              �?      @               @      �?       @               @      �?                      @      @              @       @      @              �?       @      �?                       @      >@       @      =@       @      1@      �?      @              *@      �?       @      �?              �?       @              @              (@      �?              �?      (@              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�v}hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         b                    �?��eC~�?�           8�@ �������       ]                 p�H@������?�            `n@      @       D                    �?�H�]�r�?p            @e@�aQ         	                 ��@r�0p�?F            �Z@ �aQ                             �?P���Q�?             4@       ������������������������       �        	             ,@                                ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?      @
                            @��V#�?8            �U@     �D@                           L@>A�F<�?             C@     @                           �?     ��?             @@        ������������������������       �                     @       @                        `f�)@�����H�?             ;@      �?������������������������       �                     &@      �?                           �?     ��?             0@                                  :@r�q��?             (@        ������������������������       �                      @      �?������������������������       �                     $@                                   <@      �?             @                                  �9@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @      @                        `f�2@�q�q�?             @        ������������������������       �                     @      @������������������������       �                      @      @       7                 �|�<@     ��?              H@              ,                 Ь�!@�5��?             ;@              #                   �6@���Q��?             .@               "                 �&B@�<ݚ�?             "@     �R@        !                    4@      �?             @      0@������������������������       �                      @      &@������������������������       �                      @      �?������������������������       �                     @       $       %                 �&B@�q�q�?             @      @������������������������       �                     �?     @&       '                   �9@���Q��?             @       @������������������������       �                      @      �?(       )                   �@�q�q�?             @        ������������������������       �                     �?       @*       +                 �?�@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?      ;@-       0                    �?r�q��?	             (@      @.       /                    4@�q�q�?             @      @������������������������       �                     �?       ������������������������       �                      @       @1       6                 ��.@�����H�?             "@      @2       3                   �-@z�G�z�?             @       @������������������������       �                      @        4       5                 �yG(@�q�q�?             @     �?������������������������       �                      @      �?������������������������       �                     �?       @������������������������       �                     @        8       =                 �|Y>@���N8�?             5@     �?9       :                    �?@4և���?             ,@     �?������������������������       �                     $@     "@;       <                    �?      �?             @      @������������������������       �                     �?     @������������������������       �                     @      @>       A                    @@և���X�?             @      "@?       @                    �?      �?             @      "@������������������������       �                     �?       ������������������������       �                     @      �?B       C                   �A@�q�q�?             @ 6aQ  ������������������������       �                      @ �aQ  ������������������������       �                     �? �aQ  E       J                    �?      �?*             P@      �?F       I                    �?���Q��?	             .@PaQ  G       H                 `�@1@�eP*L��?             &@       @������������������������       �                     @ "aQ  ������������������������       �                     @ "aQ  ������������������������       �                     @ (aQ  K       L                    @Rg��J��?!            �H@ �aQ  ������������������������       �                     @ �aQ  M       N                    (@��6���?             E@ -aQ  ������������������������       �                      @ �aQ  O       P                   �:@�ʻ����?             A@ aQ  ������������������������       �        
             &@        Q       \                     @�LQ�1	�?             7@aQ  R       [                    @X�<ݚ�?
             2@�aQ  S       T                   �?@��.k���?	             1@ aQ  ������������������������       �                     @�aQ  U       V                     @�q�q�?             (@ haQ  ������������������������       �                     @�LaQ  W       X                    �?      �?              @ �aQ  ������������������������       �                      @!^aQ  Y       Z                 ��p@@�q�q�?             @ aQ  ������������������������       �                     @�aQ  ������������������������       �                      @aQ  ������������������������       �                     �? aQ  ������������������������       �                     @:�aQ  ^       _                    !@��pBI�?0            @R@ aQ  ������������������������       �                     �? BaQ  `       a                    @�k~X��?/             R@�aQ  ������������������������       �        .            �Q@        ������������������������       �                     �?NaQ  c       n                    @K�(i�?"           @}@        d       i                    �?8����?             7@       e       f                     @�q�q�?             (@�aQ  ������������������������       �                     @ �aQ  g       h                 �y�-@����X�?             @ �aQ  ������������������������       �                      @ �aQ  ������������������������       �                     @^KaQ  j       k                     @"pc�
�?             &@       ������������������������       �                     @?�aQ  l       m                 pf�@@���Q��?             @ =aQ  ������������������������       �                     @aaQ  ������������������������       �                      @ aQ  o       �                    �?4�<����?           �{@ %aQ  p       {                 P�J.@����X�?4             U@ &aQ  q       r                   @@     ��?             @@�aQ  ������������������������       �                     1@ �aQ  s       z                 �(@z�G�z�?             .@        t       y                 �y�#@և���X�?             @       u       x                 �� @z�G�z�?             @       v       w                    ?@�q�q�?             @ �aQ  ������������������������       �                     �?�aQ  ������������������������       �                      @�aQ  ������������������������       �                      @ �aQ  ������������������������       �                      @        ������������������������       �                      @�aQ  |       �                    �?�E��
��?              J@aQ  }       �                   �H@j���� �?            �I@)aQ  ~       �                     @      �?             E@�aQ         �                     �?��%��?            �B@9aQ  �       �                   �8@*;L]n�?             >@ �aQ  �       �                  D�U@r�q��?             @ 910,15.������������������������       �                     �? 58,,S
6������������������������       �                     @ 0.5,,S
�       �                    �?�q�q�?             8@rgue)",�       �                 �ܵ<@      �?             4@ iss. El������������������������       �                      @,"Ander�       �                    �?r�q��?
             2@ale,39,�       �                 `f�A@      �?             (@ ,,0,0,S������������������������       �                     @  Jane",�       �                 @�6M@      �?             @ e,,0,0,������������������������       �                     @ male,35������������������������       �                     @ 24,1,2,������������������������       �                     @ 1,1,347�       �                 @��v@      �?             @K Stanl������������������������       �                     @ss. Mar������������������������       �                     �? r. Lawr������������������������       �                     @ oni",ma�       �                    �?z�G�z�?             @ son Jr"������������������������       �                     �?id",male������������������������       �                     @ard",ma������������������������       �                     "@  ""Dai"������������������������       �                     �?ick",mal�       �                 `ff:@���5���?�            �v@les Leo�       �                    �?��S�jC�?�            pr@ Gretch�       �                    )@(�s���?�            �o@ ndyeff,������������������������       �                      @nnell, �       �                   @E@ ��GS=�?�            @o@rth, Mr�       �                   �D@�IєX�?�            �k@,3,"Lun�       �                 ���@�X�<ݺ?�             k@ 3,1,1,"������������������������       �                    �C@ 34,0,1,�       �                 �?$@ ,��-�?i             f@ ,0,3,"S�       �                   �;@�㙢�c�?             7@ avis, M������������������������       �                     @ Mr. Ant�       �                    �?������?
             1@,"Colly�       �                 �|Y=@d}h���?             ,@ Panula,������������������������       �                      @ .6875,,������������������������       ��8��8��?             (@6.1,,S
�       �                 �|Y?@�q�q�?             @ 2,,S
64������������������������       �                     �? B35,C
6������������������������       �                      @ 8,27.9,�       �                 �?�@�kb97�?[            @c@ 5,1,3,"������������������������       �                    �A@ 46,1,1,�       �                   �3@T(y2��?C            �]@ D33,C
6�       �                   �1@��2(&�?             6@ 48,1,1,������������������������       �                     @35.5,A26�       �                 0S5 @z�G�z�?	             .@ .55,,S
�       �                   �2@      �?             @ A. 2314������������������������       �                     �?958,,S
������������������������       ��q�q�?             @ 653,0,3������������������������       �                     &@,,S
654�       �                    �?h�a��?7            @X@,7.8292�       �                 �|�=@ rpa�?5            @W@0,36522�       �                 @3�!@��v$���?!            �N@ ,S.O.C.�       �                 pf� @�nkK�?             7@349223,������������������������       �        
             4@32,1,1,�       �                    8@�q�q�?             @ e,23,0,������������������������       �                      @8,0,2,3������������������������       �                     �? ",male,������������������������       �                     C@e,40,0,�       �                   �?@      �?             @@ ,47,0,0�       �                     @�<ݚ�?             "@ 0,34921������������������������       �                     @,1,0,ST�       �                 @3�@      �?             @ e,32,2,������������������������       �                     �?on",mal�       �                 �̌!@�q�q�?             @ ",male,������������������������       �                      @ 0,A/5 3������������������������       �                     �?ummins W�       �                   �@@���}<S�?             7@ Thomas ������������������������       �                     "@ ,29750,�       �                     @؇���X�?	             ,@2750,52�       �                   �3@؇���X�?             @C.A. 24�       �                   �A@r�q��?             @ 44270,1������������������������       ��q�q�?             @ 6,0,,S
������������������������       �                     @12,7.77������������������������       �                     �? 0,34282�       �                 @3�@؇���X�?             @ ,4138,9������������������������       ��q�q�?             @",femal������������������������       �                     @ ke Mart������������������������       �                     @ ,"Peter�       �                 ���%@z�G�z�?             @ sab, Mr������������������������       �                     @ vigen, ������������������������       �      �?              @dwin, M������������������������       �                     =@ rown, M�       �                     @ qP��B�?            �E@ 2,"Laro������������������������       �                      @ 2123,41�       �                   �/@��?^�k�?            �A@101295,������������������������       �                     2@,10.170�       �                    )@�IєX�?             1@ 0,35003������������������������       �                     �? emale,1������������������������       �        
             0@ n",male�       �                    �?:ɨ��?-            �P@e,4,0,1�       �                    �?���Q��?              I@56.4958�       �                     �?��.k���?             A@695,0,1�       �                   �>@X�<ݚ�?             ;@hapman,�       �                    R@����X�?             5@elly, M�       �                   @=@�q�q�?             2@ss. Kat�       �                 �|�<@���Q��?             $@ ayer, M������������������������       �                     �?,"Humbl�       �                 `f�;@�q�q�?             "@.65,F G�       �                 �|�?@      �?              @ Force)"������������������������       �                     @thorne,�       �                   �J@���Q��?             @ 03,0,3,������������������������       �                     @,0,3,"G������������������������       �                      @,"Hanse������������������������       �                     �?"Morley������������������������       �                      @ 50655,2������������������������       �                     @ 0,0,223������������������������       �                     @male,42,�       �                 �|�>@؇���X�?             @,female������������������������       �                     @  Gonios������������������������       �                     �?,"Mayne,�       �                 ��9L@      �?
             0@,0,PC 1�       �                   �C@ףp=
�?             $@ ,113028������������������������       �                     @1,0,199�       �                    G@�q�q�?             @,0,0,75�       �                     �?      �?              @ 250647,������������������������       �                     �? ",male,������������������������       �                     �?e Louis������������������������       �                     �? Miss. E�       �                   �D@      �?             @19,0,3,�       �                     �?      �?             @hnson, ������������������������       �                     @,"Harper������������������������       �                     �?722,0,3������������������������       �                      @
723,0,������������������������       �                     0@724,0,2�t�b��     h�h*h-K ��h/��R�(KK�KK��h]�B�       p|@      p@     �O@     �f@     �N@     @[@      =@     @S@      �?      3@              ,@      �?      @              @      �?              <@      M@      @      ?@      @      =@              @      @      8@              &@      @      *@       @      $@       @                      $@      �?      @      �?      �?              �?      �?                       @      @       @      @                       @      5@      ;@      0@      &@      @      "@       @      @       @       @       @                       @              @      @       @      �?              @       @       @              �?       @              �?      �?      �?      �?                      �?      $@       @       @      �?              �?       @               @      �?      @      �?       @               @      �?       @                      �?      @              @      0@      �?      *@              $@      �?      @      �?                      @      @      @      @      �?              �?      @              �?       @               @      �?              @@      @@      "@      @      @      @      @                      @      @              7@      :@              @      7@      3@       @              .@      3@              &@      .@       @      $@       @      "@       @      @              @       @              @      @      @       @               @      @              @       @              �?              @               @     �Q@      �?              �?     �Q@             �Q@      �?             �x@      S@      @      0@      @      @              @      @       @               @      @               @      "@              @       @      @              @       @             x@      N@      N@      8@      =@      @      1@              (@      @      @      @      @      �?       @      �?              �?       @               @                       @       @              ?@      5@      >@      5@      5@      5@      4@      1@      *@      1@      @      �?              �?      @               @      0@      @      .@       @              @      .@      @      "@              @      @      @      @                      @              @      @      �?      @                      �?      @              �?      @      �?                      @      "@              �?             Pt@      B@     pq@      0@     �m@      .@               @     �m@      *@      j@      *@     �i@      (@     �C@             �d@      (@      3@      @      @              *@      @      &@      @               @      &@      �?       @      �?              �?       @             @b@       @     �A@             �[@       @      3@      @      @              (@      @      �?      @              �?      �?       @      &@              W@      @      V@      @      N@      �?      6@      �?      4@               @      �?       @                      �?      C@              <@      @      @       @      @               @       @              �?       @      �?       @                      �?      5@       @      "@              (@       @      @      �?      @      �?       @      �?      @              �?              @      �?       @      �?      @              @              @      �?      @              �?      �?      =@              E@      �?       @              A@      �?      2@              0@      �?              �?      0@              G@      4@      >@      4@      2@      0@      (@      .@      @      .@      @      (@      @      @              �?      @      @      @      @      @               @      @              @       @              �?                       @              @      @              @      �?      @                      �?      (@      @      "@      �?      @               @      �?      �?      �?              �?      �?              �?              @      @      �?      @              @      �?               @              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg}�XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMChuh*h-K ��h/��R�(KMC��h|�B�P         r                 `f�$@��t���?�           8�@      G@                            @z�G�z�?�            @p@        ������������������������       �                      @     @       k                   @@@Z���c��?�            �o@�aQ                              �?�۲I <�?�            �j@                                �|Y=@T�7�s��?#            �L@                                ���@"pc�
�?             &@               	                   �2@�q�q�?             @        ������������������������       �                     �?���XQ  
                        �{@      �?              @ ��XQ  ������������������������       �                     �?���XQ  ������������������������       �                     �?ppDYQ  ������������������������       �                      @���XQ                          03@�LQ�1	�?             G@\�XQ                          ���@���"͏�?            �B@ ��XQ                             �?$�q-�?             *@ ��XQ  ������������������������       �                     �?      @������������������������       �                     (@      @                           �?�q�q�?             8@     @                        ��@�LQ�1	�?             7@       @������������������������       �                      @       @                           �?����X�?             5@     @                           �?�q�q�?             2@      @������������������������       �                     @       @                        ���@؇���X�?	             ,@       @������������������������       �                     �?        ������������������������       �8�Z$���?             *@        ������������������������       �                     @     @U@������������������������       �                     �?                                   �?�<ݚ�?             "@    �I@������������������������       �                     @      &@������������������������       �                      @        !       4                    �?�IA��?e            �c@      @"       3                 �|Y>@     ��?             0@       #       2                    �?���Q��?             .@     6@$       -                   �6@և���X�?             ,@     ,@%       ,                 xF� @X�<ݚ�?             "@     @&       +                    �?r�q��?             @     �?'       *                   �3@z�G�z�?             @        (       )                 P��@      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      >@������������������������       �                     @      �?������������������������       �                     �?        ������������������������       �                     @       @.       /                 �&B@z�G�z�?             @      @������������������������       �                      @       @0       1                    9@�q�q�?             @     �?������������������������       �                      @      �?������������������������       �                     �?      �?������������������������       �                     �?      @������������������������       �                     �?      @5       H                 �?�@`	�<��?V            �a@     �?6       E                   �?@��p\�?.            �T@     �?7       <                 ���@ �\���?,            �S@        8       9                    7@����X�?             @        ������������������������       �                     @        :       ;                 �&b@      �?             @     @������������������������       �                      @      H@������������������������       �                      @      @=       D                 �?$@������?'             R@        >       ?                 �|Y;@HP�s��?             9@       ������������������������       �        
             2@      �?@       C                 �|Y>@����X�?             @     7@A       B                 ��@���Q��?             @      @������������������������       �                     @      �?������������������������       �                      @      �?������������������������       �                      @        ������������������������       �                    �G@        F       G                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       R                 @3�@��$�4��?(            �M@        J       Q                    �?X�<ݚ�?             "@       K       P                    �?      �?              @       L       M                   �9@և���X�?             @        ������������������������       �                      @        N       O                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        S       h                 �|�=@j�q����?"             I@       T       a                 @�!@��0{9�?             �G@       U       ^                   � @"pc�
�?            �@@       V       ]                 0S5 @�>4և��?             <@       W       \                   �4@�+$�jP�?             ;@        X       Y                    1@X�<ݚ�?             "@        ������������������������       �      �?             @        Z       [                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     2@        ������������������������       �                     �?        _       `                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        b       c                 ���"@@4և���?
             ,@        ������������������������       �                     @        d       e                   �<@ףp=
�?             $@       ������������������������       �                     @        f       g                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        i       j                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        l       m                   @C@P�Lt�<�?             C@        ������������������������       �                     3@        n       o                    �?�}�+r��?             3@        ������������������������       �                      @        p       q                   �C@�IєX�?
             1@        ������������������������       ��q�q�?             @        ������������������������       �                     ,@        s                           @.iI\��?           0|@       t       �                  x#J@$;hB��?�            @s@       u       �                   �<@��U��?�            �j@        v       �                    �?��V#�?1            �U@       w       x                    �?@3����?             K@        ������������������������       �                      @        y       �                    �?��<b�ƥ?             G@        z       {                   �6@�nkK�?	             7@        ������������������������       �                     "@        |                          �9@@4և���?             ,@        }       ~                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     7@        �       �                    �?     ��?             @@        �       �                    �?և���X�?             @       �       �                   �8@���Q��?             @       �       �                 hf:@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@HP�s��?             9@       ������������������������       �                     7@        ������������������������       �                      @        �       �                    �?b����?R            �_@       �       �                  �?@�8�Վ��?Q            @_@       �       �                    �?D��ٝ�?B            @Y@        �       �                    �?�eP*L��?             6@        �       �                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?       �       �                   @C@     ��?	             0@       �       �                 ��";@r�q��?             (@       �       �                   @@@�q�q�?             @        ������������������������       �                     @        �       �                   �A@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                     @       �       �                     �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���%&�?5            �S@       �       �                   �F@^H���+�?2            �R@       �       �                   @F@�[�IJ�?             �G@       �       �                   @E@�lg����?            �E@       �       �                     �?�e����?            �C@        �       �                 �|�?@�q�q�?             @       �       �                   �>@z�G�z�?             @       �       �                 `f�;@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �C@4���C�?            �@@       �       �                   @B@����"�?             =@       �       �                    �?
;&����?             7@        ������������������������       �                     "@        �       �                    1@؇���X�?             ,@       �       �                   �'@�<ݚ�?             "@        ������������������������       �                     @       �       �                    @@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @       �       �                   �,@      �?             @        ������������������������       �      �?              @       ������������������������       �                      @        ������������������������       �                     @       ������������������������       �                     @        �       �                   �R@�<ݚ�?             ;@       �       �                    �?���B���?             :@        ������������������������       �                     @        �       �                    �?���}<S�?             7@       �       �                   �I@�C��2(�?             6@       �       �                 ��:@r�q��?             (@       ������������������������       �                      @        �       �                 `f�;@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@       ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             8@        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                     �?        �                         �O@�q�q�?A             X@       �       �                   �5@���!pc�?>             V@        �       �                   �1@��.k���?             1@       �       �                 ��f`@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       �       �                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @       �       �                 `fmj@@���?T�?3            �Q@       �       �                    �?     8�?.             P@       �       �                 ���P@���-T��?-             O@        �       �                 03sP@�z�G��?             4@       �       �                    �?@�0�!��?             1@        ������������������������       �                     $@        �       �                   �H@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                 0�nL@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @        ������������������������       �                     @        �       �                    �?@4և���?              E@       �       �                    �?@-�_ .�?            �B@       �       �                    �?`Jj��?             ?@       ������������������������       �                     0@       �       �                    �?�r����?             .@        ������������������������       �                     @       �       �                   �H@      �?              @       �       �                 ЈT@؇���X�?             @        ������������������������       �                     @       �       �                   �D@      �?             @        ������������������������       �                      @        �       �                 Ј�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��W@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?և���X�?             @        ������������������������       �                     �?       �                          �?      �?             @                              �̾w@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                 �?x�f��^�?[            �a@                                 �?�>$�*��?            �D@                             X�,A@��+7��?             7@             	                  �0@��s����?             5@        ������������������������       �                     @        
                        �7@������?             .@        ������������������������       �                     �?                              �|Y=@d}h���?             ,@        ������������������������       �                      @                                 �?      �?             (@                              S�-@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             2@                             03�-@�eP*L��?             &@                                 3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r�q��?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              8                   �?t�F�}�?B            �Y@              /                   �?�q�q�?'             N@        !      *                ���5@*;L]n�?             >@       "      )                  �D@     ��?
             0@       #      (                   7@�r����?	             .@        $      '                   �?      �?             @       %      &                   +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        +      .                  @C@����X�?             ,@        ,      -                X��@@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0      1                   )@������?             >@        ������������������������       �                     @        2      7                   ;@H%u��?             9@        3      6                   �?և���X�?             @        4      5                �!&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        9      B                   @@4և���?             E@        :      ;                   �?���!pc�?             &@        ������������������������       �                     @        <      =                   @և���X�?             @        ������������������������       �                     @        >      ?                   �?      �?             @        ������������������������       �                      @        @      A                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �t�bh�h*h-K ��h/��R�(KMCKK��h]�B0       �{@     �p@      j@      J@       @              i@      J@     `d@     �I@      @@      9@       @      "@       @      �?      �?              �?      �?      �?                      �?               @      >@      0@      <@      "@      (@      �?              �?      (@              0@       @      .@       @               @      .@      @      (@      @              @      (@       @      �?              &@       @      @              �?               @      @              @       @             ``@      :@      "@      @      "@      @       @      @      @      @      �?      @      �?      @      �?      �?              �?      �?                      @              �?      @              @      �?       @               @      �?       @                      �?      �?                      �?     �^@      3@      S@      @     �R@      @      @       @      @               @       @       @                       @     �Q@       @      7@       @      2@              @       @      @       @      @                       @       @             �G@              �?       @               @      �?              G@      *@      @      @      @      @      @      @       @               @      @              �?       @       @              �?      �?             �D@      "@      D@      @      ;@      @      7@      @      6@      @      @      @      @      �?      �?      @               @      �?       @      2@              �?              @      �?      @                      �?      *@      �?      @              "@      �?      @               @      �?              �?       @              �?       @               @      �?             �B@      �?      3@              2@      �?       @              0@      �?       @      �?      ,@             @m@      k@     �a@     �d@     �[@     �Y@      <@      M@      �?     �J@               @      �?     �F@      �?      6@              "@      �?      *@      �?      @      �?                      @              "@              7@      ;@      @      @      @       @      @       @      �?       @                      �?               @       @              7@       @      7@                       @     �T@      F@     �T@     �E@     �N@      D@      (@      $@      �?      @              @      �?              &@      @      $@       @      @       @      @              �?       @               @      �?              @              �?      @              @      �?             �H@      >@      H@      :@      ;@      4@      ;@      0@      7@      0@      @       @      @      �?      �?      �?      �?                      �?      @                      �?      3@      ,@      2@      &@      (@      &@              "@      (@       @      @       @      @              @       @      @              �?       @      @              @              �?      @      �?      �?               @      @                      @      5@      @      5@      @              @      5@       @      4@       @      $@       @       @               @       @               @       @              $@              �?                      �?      �?      @      �?                      @      5@      @              @      5@                      �?      @@      P@      8@      P@      "@       @      �?      @              @      �?      �?      �?                      �?       @       @       @                       @      .@      L@      &@     �J@      "@     �J@      @      ,@      @      ,@              $@      @      @      �?      @              @      �?      �?              �?      �?               @              @              @     �C@       @     �A@       @      =@              0@       @      *@              @       @      @      �?      @              @      �?      @               @      �?      �?      �?                      �?      �?                      @      �?      @              @      �?               @              @      @      �?              @      @      @       @      @                       @              �?       @              W@     �I@      2@      7@      @      1@      @      1@              @      @      &@      �?              @      &@               @      @      "@      @      @      @                      @               @       @              (@      @      @      @      @      �?              �?      @              �?      @      �?      �?      �?                      �?              @      @             �R@      <@     �A@      9@      *@      1@      @      *@       @      *@       @       @       @      �?              �?       @                      �?              &@      �?              $@      @      @      @      @                      @      @              6@       @              @      6@      @      @      @      �?      @      �?                      @      @              2@             �C@      @       @      @      @              @      @      @              �?      @               @      �?      �?      �?                      �?      ?@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ	�tlhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         J                    �?�4�O��?�           8�@               5                    �?r�=���?~            �h@                                  �?T �����?[             c@      =@                           �?�i�y�?$            �O@     *@                           �?`Ӹ����?            �F@        ������������������������       �                     6@      3@                            @���}<S�?             7@      *@������������������������       �                     @      &@	       
                 ���@�����H�?             2@       ������������������������       �                      @       ������������������������       �        
             0@       ������������������������       �        
             2@                                    �?��Hg���?7            �V@                                   �?և���X�?             5@                                  �?���Q��?             4@                               `f�A@�q�q�?             (@      ������������������������       �                     @      @������������������������       �                     @      @                          �5@      �?              @      @������������������������       �                      @       @                          �H@r�q��?             @      @������������������������       �                     @     @������������������������       �                     �?      @������������������������       �                     �?       @                        ���@�~t��?*            @Q@       @������������������������       �        
             2@               4                    �?��x_F-�?             �I@              3                 �|�=@j�q����?             I@    @U@       *                    �?      �?             B@              %                   �:@���y4F�?             3@     �I@                         �&�)@�q�q�?             @      &@������������������������       �                     �?        !       "                   �8@z�G�z�?             @      �?������������������������       �                     @     8@#       $                 �0@      �?              @        ������������������������       �                     �?      4@������������������������       �                     �?      &@&       )                   @@8�Z$���?             *@        '       (                 �|=@�q�q�?             @        ������������������������       �                      @      �?������������������������       �      �?             @      @������������������������       �                     @      @+       .                 �|Y=@�t����?
             1@      �?,       -                  ��@      �?             @      �?������������������������       �                      @      �?������������������������       �                      @      @/       2                    �?�θ�?             *@     �?0       1                  s�@�z�G��?             $@      �?������������������������       �                     @        ������������������������       �      �?             @       @������������������������       �                     @      @������������������������       �                     ,@      @������������������������       �                     �?       @6       C                    �?8�A�0��?#             F@     @7       <                 �|Y=@�LQ�1	�?             7@     �?8       ;                 03�-@r�q��?
             (@      $@9       :                    &@�q�q�?             @      @������������������������       �                     �?      @������������������������       �                      @       @������������������������       �                     "@        =       B                    �?�eP*L��?	             &@       >       ?                   @E@r�q��?             @        ������������������������       �                     @      �?@       A                 <3gH@�q�q�?             @       @������������������������       �                     �?        ������������������������       �                      @      1@������������������������       �                     @      &@D       I                     @؇���X�?             5@       E       H                 �̾w@�θ�?             *@     @F       G                    )@�C��2(�?
             &@        ������������������������       �                     �?      �?������������������������       �        	             $@      9@������������������������       �                      @       @������������������������       �                      @      �?K       �                    �?D����?C           �@      @L       m                    �?�BA����?f            `d@       @M       l                   �J@�7�QJW�?/            �R@     @N       [                     @v���a�?.            @R@       O       P                   �6@$�q-�?             J@      @������������������������       �        	             2@      �?Q       Z                   �*@�t����?             A@        R       S                   �'@�	j*D�?
             *@        ������������������������       �                      @        T       U                    :@���|���?             &@        ������������������������       �                      @        V       W                   �B@�<ݚ�?             "@       ������������������������       �                     @        X       Y                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        \       k                    @�q�q�?             5@       ]       j                 @�"@�z�G��?             4@       ^       i                 `��!@և���X�?
             ,@       _       b                 ���@�q�q�?	             (@        `       a                 �|Y:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        c       d                    4@և���X�?             @        ������������������������       �                      @        e       f                 @3�@z�G�z�?             @       ������������������������       �                     @        g       h                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        n       �                 �D�H@��7��?7             V@       o       �                    @�{r٣��?'            �P@       p       q                    @JJ����?            �G@        ������������������������       �                     @        r       �                    �?�D����?             E@       s       �                    @\�Uo��?             C@       t       u                   �6@և���X�?            �A@        ������������������������       �                     @        v       }                     @     ��?             @@        w       x                   �7@      �?             (@        ������������������������       �                      @        y       |                    �?ףp=
�?             $@       z       {                    D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~                        �|Y=@�z�G��?             4@        ������������������������       �                     @        �       �                    �?���Q��?             .@        �       �                 ��1@�q�q�?             @,0,SOTO������������������������       �                     @ ,,1,0,3������������������������       �                      @ le,30,0�       �                 `fV6@�<ݚ�?             "@ a Sophi������������������������       �                     �? ussa, M�       �                 ��T?@      �?              @,"Jermy������������������������       �                     @t, Mme. ������������������������       �                     �?1,1,"Har������������������������       �                     @C
372,0,�       �                    �?      �?             @ ,S
373,������������������������       �                      @,,S
374,������������������������       �                      @,C
375,0�       �                 pfv2@p�ݯ��?
             3@ 5,,S
37������������������������       �                     @ ,PC 176�       �                    �?$�q-�?             *@ emale,2������������������������       �                      @ male,27�       �                 ��T?@z�G�z�?             @e,20,0,������������������������       �                     @ale,19,0������������������������       �                     �?e,42,0,0�       �                    #@�C��2(�?             6@ ")",fem������������������������       �                     �?ale,32,0�       �                 ���P@���N8�?             5@ exander������������������������       �                     $@ 5,0,3,"�       �                 X�,@@�C��2(�?             &@ 2,"Davi�       �                    �?�q�q�?             @ 87,0,3,������������������������       �                     �?,,S
388�       �                 ���d@      �?              @ ,"Sadli������������������������       �                     �?mann, Mi������������������������       �                     �? Mr. Wil������������������������       �                      @ nsson, �       �                     �?PN��T'�?�            �u@ afsson,�       �                   �>@�j�'�=�?*            �P@ Newell,�       �                   �<@r�q��?             8@ 3,"Sand������������������������       �                     @4,0,2,P�       �                   �Q@��Q��?             4@0,35005�       �                   @E@�E��ӭ�?             2@50407,7�       �                 03:@d}h���?
             ,@ 403,26,������������������������       �                      @400,1,2�       �                 03k:@      �?             @ 12.65,,������������������������       �                     �? 289,7.9�       �                 �|�?@���Q��?             @S
403,0�       �                 `fF<@      �?             @ 
404,0,������������������������       �                      @3101279,�       �                 �|Y=@      �?              @ 315096,������������������������       �                     �?,21,,S
4������������������������       �                     �? 064,7.7������������������������       �                     �?,29106,1�       �                    K@      �?             @21,0,0,�       �                   @G@�q�q�?             @4133,25������������������������       �      �?              @.8958,,S������������������������       �                     �?3,1,1,"M������������������������       �                     �?0,2,"Cun������������������������       �                      @ 3,"Sund�       �                 �|�<@��s����?             E@ 5,,S
41������������������������       �                     @0,0,3430�       �                    �?�ݜ�?            �C@Christi�       �                   �E@4?,R��?             B@yyli Ka�       �                  x#J@�E��ӭ�?             2@. Willi������������������������       �                     "@. Cathar�       �                 �|Y>@X�<ݚ�?             "@ r. Stan������������������������       �                      @ id",mal�       �                 `f�K@����X�?             @ ",male,�       �                 `�iJ@�q�q�?             @ t (Anna������������������������       �                     �?0,3,"Ro������������������������       �                      @426,0,3������������������������       �                     @ 7,1,2,"������������������������       �        	             2@,0,2003,������������������������       �                     @ Louise �       �                    '@�W�{�5�?�            �q@ "Flynn,�       �                     @��H�}�?             9@ . Berk ������������������������       �                     @,S
431,1�       �                 ���A@      �?
             2@0,11056�       �                    @ףp=
�?             $@ nce Kat������������������������       �                     �? Charle������������������������       �                     "@085,26,,������������������������       �                      @O 2. 310�       �                 �?�@0Oex�I�?�            @p@ ,1,0,13�       �                     @p� V�?=            �Y@ ,14,1,2������������������������       �                     @ et ""Da�       �                    ?@@��8��?9             X@ds, Mrs�       �                   �8@@�z�G�?.             T@ 9,0,1,"�       �                    7@ ���J��?            �C@0,0,2,"������������������������       �                     ?@ 18723,1�       �                 `fF@      �?              @ d)",fem�       �                 �&b@�q�q�?             @ ",male,������������������������       �                      @,male,25������������������������       �                     �?female,������������������������       �                     @ Bernt",������������������������       �                    �D@ ton",ma�       �                 �&B@      �?             0@deleine������������������������       �        
             .@r. Frede������������������������       �                     �? Miss. �                          �?P��-�?h            �c@uchen, �       �                     @0�I��8�?T             _@ ,0,2,"W�       �                    F@dP-���?!            �G@,0,3,"H�       �                   @D@������?            �B@S
453,0�       �                   �3@�#-���?            �A@7.75,C1�       �                   �(@ȵHPS!�?             :@ ,89.104�       �                   �5@$�q-�?             *@ 8.05,,S�       �                    &@r�q��?             @ C
457,0������������������������       �                     �?38,S
458������������������������       �                     @64,51.86������������������������       �                     @C. 1353�       �                 �|�<@8�Z$���?
             *@ 0,7.75,������������������������       �                     @E12,S
4�       �                   �A@�q�q�?             @63,0,1,�       �                 �|�=@�q�q�?             @ ,"Milli������������������������       �                     �?3,"Maisn�       �                    @@      �?              @ ves, Mr������������������������       �                     �?,S
467,0������������������������       �                     �?,"Smart,������������������������       �                     @ ,"Scanl������������������������       �                     "@ Miss. ������������������������       �      �?              @Keefe, ������������������������       �                     $@Luka",m�                         @@@؇���X�?3            @S@ur (Ada�       
                �|Y>@���*�?&             N@Jerwan,�                       �!&B@�t����?!            �I@H Basle�       �                   �1@�8��8��?             H@ male,22������������������������       �                     $@",male,,�       �                   �2@�KM�]�?             C@ e,34,1,������������������������       �                     �?9,1,0,34�       �                 ��) @�L���?            �B@ 0,0,350������������������������       �                     4@,0,1,31�                       @3�!@@�0�!��?             1@ ,male,9�       �                 pf� @�q�q�?             @ rchie""������������������������       �                     �?y",male,                       �|Y<@      �?              @ female,������������������������       �                     �?       ������������������������       �                     �?                               �<@@4և���?             ,@       ������������������������       �                     &@                             �|Y=@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @             	                   ;@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?                               �?@X�<ݚ�?             "@ � 6�t� ������������������������       �                     @                              ��I @�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                    �@@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B       �{@     �p@      X@     @Y@     �Q@     �T@       @     �N@       @     �E@              6@       @      5@              @       @      0@       @                      0@              2@      Q@      6@      "@      (@       @      (@      @      @              @      @              @      @       @              �?      @              @      �?              �?             �M@      $@      2@             �D@      $@     �D@      "@      ;@      "@      .@      @      @       @              �?      @      �?      @              �?      �?      �?                      �?      &@       @      @       @       @               @       @      @              (@      @       @       @       @                       @      $@      @      @      @      @              @      @      @              ,@                      �?      :@      2@       @      .@       @      $@       @      �?              �?       @                      "@      @      @      �?      @              @      �?       @      �?                       @      @              2@      @      $@      @      $@      �?              �?      $@                       @       @             �u@     `d@      J@     �[@      *@      O@      &@      O@      @      H@              2@      @      >@      @      "@               @      @      @       @               @      @              @       @      �?       @                      �?              5@      @      ,@      @      ,@      @       @      @       @      �?      @              @      �?              @      @       @              �?      @              @      �?      �?      �?                      �?       @                      @      �?               @             �C@     �H@     �B@      =@      9@      6@              @      9@      1@      7@      .@      4@      .@      @              1@      .@      @      "@       @              �?      "@      �?      @              @      �?                      @      ,@      @      @              "@      @       @      @              @       @              @       @              �?      @      �?      @                      �?      @               @       @               @       @              (@      @              @      (@      �?       @              @      �?      @                      �?       @      4@      �?              �?      4@              $@      �?      $@      �?       @              �?      �?      �?      �?                      �?               @     �r@      J@     �G@      3@      *@      &@              @      *@      @      *@      @      &@      @       @              @      @              �?      @       @      @      �?       @              �?      �?      �?                      �?              �?       @       @      �?       @      �?      �?              �?      �?                       @      A@       @              @      A@      @      ?@      @      *@      @      "@              @      @       @               @      @       @      �?              �?       @                      @      2@              @             �o@     �@@      "@      0@              @      "@      "@      �?      "@      �?                      "@       @             `n@      1@     @Y@       @      @             �W@       @     �S@      �?      C@      �?      ?@              @      �?       @      �?       @                      �?      @             �D@              .@      �?      .@                      �?     �a@      .@     @[@      .@     �E@      @     �@@      @      @@      @      7@      @      (@      �?      @      �?              �?      @              @              &@       @      @              @       @      �?       @              �?      �?      �?      �?                      �?      @              "@              �?      �?      $@             �P@      &@     �H@      &@     �F@      @      F@      @      $@              A@      @              �?      A@      @      4@              ,@      @      �?       @              �?      �?      �?              �?      �?              *@      �?      &@               @      �?              �?       @              �?       @               @      �?              @      @              @      @       @      @       @      �?              1@             �@@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ޡhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         �                 `f~I@�t����?�           8�@              S                    �?�����2�?�           h�@      �?                        ��@V���#�?~            �g@      2@                        �|Y:@�IєX�?             1@     @������������������������       �                     &@��aQ                          �&�@r�q��?             @      3@������������������������       �                     �?     @������������������������       �                     @4�aQ  	                            @�.�8�?q            �e@        
                        ���*@�L#���?/            �P@                                `f�)@      �?             8@                                  �J@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?                                 �B@"pc�
�?	             &@                                  :@�����H�?             "@                                   �?�q�q�?             @      @������������������������       �                     �?        ������������������������       �                      @     �[@������������������������       �                     @      2@                           D@      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      ,@                           E@ qP��B�?            �E@     @������������������������       �                     ?@                                    �?�8��8��?             (@        ������������������������       �                     @                                   �?r�q��?             @      6@������������������������       �                     �?      .@������������������������       �                     @               &                    @�k��V��?B            �Z@                %                    �?؇���X�?             ,@     @!       $                    @      �?              @      0@"       #                 ��0@      �?             @      "@������������������������       �                      @      @������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     @      0@'       D                 03�1@�+Fi��?;             W@     *@(       =                 �?�-@�ݜ����?'            �M@     @)       ,                 �̌@�&!��?            �E@       @*       +                   �2@�z�G��?             $@        ������������������������       �                     @      @������������������������       �                     @      �?-       .                   �1@:ɨ��?            �@@      @������������������������       �                     @      �?/       <                    �?PN��T'�?             ;@     @0       1                 `�X!@���y4F�?             3@      �?������������������������       �                     @       @2       7                   �9@����X�?	             ,@     �?3       6                    4@      �?              @      �?4       5                    �?�q�q�?             @      �?������������������������       �                      @      �?������������������������       �                     �?      �?������������������������       �                     @      4@8       9                    �?      �?             @      (@������������������������       �                     �?      @:       ;                    A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @      @������������������������       �                      @      �?>       ?                   �0@      �?
             0@      @������������������������       �                     �?        @       C                   �;@��S�ۿ?	             .@        A       B                    �?�q�q�?             @        ������������������������       �                     �?       @������������������������       �                      @      @������������������������       �                     (@        E       H                    @"pc�
�?            �@@       F       G                    �?�����?             5@        ������������������������       �                      @        ������������������������       �                     3@        I       J                 0C�7@�q�q�?             (@        ������������������������       �                     �?        K       L                    �?���!pc�?             &@        ������������������������       �                     @        M       N                    @      �?              @        ������������������������       �                      @        O       R                    @      �?             @       P       Q                   @C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        T       m                 �?�@б΅t�?           �x@        U       l                    �?�wY;��?X             a@       V       k                 �Yu@     x�?S             `@       W       b                    �?���F6��?B            �X@        X       Y                 ���@�ݜ�?            �C@        ������������������������       �        	             .@        Z       [                   �6@�q�q�?             8@        ������������������������       �                      @        \       ]                  ��@��2(&�?             6@        ������������������������       �                     "@        ^       _                 �|Y=@�θ�?	             *@        ������������������������       �                     �?        `       a                 X��A@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        c       d                    7@(;L]n�?)             N@        ������������������������       �                     3@        e       j                 ��L@������?            �D@       f       g                 ���@�(\����?             D@        ������������������������       �                     5@        h       i                 ���@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                      @        n       �                     �?|;�c� �?�            pp@        o       t                 �|�<@�q�q�?              H@        p       q                   �;@؇���X�?             @        ������������������������       �                      @        r       s                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        u       �                    �?���?            �D@       v       �                  �>@�d�����?             C@       w       �                    K@���Q��?             9@       x       �                   �G@���Q��?
             .@       y       ~                    �?���Q��?             $@        z       {                 `f&;@      �?             @        ������������������������       �                      @        |       }                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                 03k:@      �?             @        �       �                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?  aQ  ������������������������       �                      @0aQ  ������������������������       �                     @ �aQ  �       �                 ���=@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @ aQ  �       �                    �?��ݼ��?�            �j@�aQ  �       �                     @�r����?W            �`@        �       �                    �? "��u�?              I@ �aQ  ������������������������       �                     �?       �       �                    �?��<D�m�?            �H@       �       �                   �*@      �?             H@       �       �                 `fF)@l��\��?             A@        ������������������������       �                     $@ ,aQ  �       �                 �|�<@      �?             8@        ������������������������       �                     *@       �       �                   �F@���!pc�?             &@       �       �                 �|�=@      �?             @ �aQ  ������������������������       �                     �? vaQ  �       �                    B@���Q��?             @        ������������������������       �                      @ aQ  ������������������������       ��q�q�?             @        ������������������������       �                     @�aQ  ������������������������       �                     ,@        ������������������������       �                     �? |aQ  �       �                    �?@�0�!��?7            @U@        ������������������������       �                     @        �       �                 @3�@����!�?4            �T@ kaQ  �       �                    :@�eP*L��?             &@        ������������������������       �                     @        �       �                   �?@����X�?             @ �aQ  ������������������������       �                      @       �       �                   �A@���Q��?             @        ������������������������       ��q�q�?             @       ������������������������       �      �?              @ �aQ  �       �                    )@D��\��?-            �Q@        ������������������������       �                     �?        �       �                 �|Y=@������?,            �Q@        �       �                 ��Y @��a�n`�?             ?@ ?aQ  �       �                   �3@      �?              @        ������������������������       �                     @�aQ  ������������������������       �                     @        �       �                 `�X#@�㙢�c�?             7@	aQ  �       �                 ���"@���y4F�?             3@FaQ  �       �                 @�!@�r����?
             .@       �       �                 pf� @�<ݚ�?             "@        ������������������������       �                      @ �aQ  �       �                    8@����X�?             @?aQ  ������������������������       �                     @ �aQ  ������������������������       �                      @        ������������������������       �                     @'aQ  �       �                   �<@      �?             @       ������������������������       �                      @saQ  ������������������������       �                      @        ������������������������       �                     @ �aQ  �       �                   �?@�7��?            �C@�aQ  �       �                 ��) @���}<S�?             7@       ������������������������       �                     ,@	aQ  �       �                 �|�=@�<ݚ�?             "@aQ  �       �                 pf� @      �?              @ �aQ  ������������������������       �                     �? �aQ  ������������������������       �                     @       ������������������������       �                     �?       ������������������������       �        	             0@ �aQ  �       �                    �?�z�G��?5             T@ �aQ  �       �                 �2@�n_Y�K�?             *@       �       �                 �|�;@�����H�?             "@       �       �                 �&�)@      �?             @ �aQ  ������������������������       �                      @ DaQ  �       �                    �?      �?              @ aQ  ������������������������       �                     �?        ������������������������       �                     �? �aQ  ������������������������       �                     @        ������������������������       �                     @3aQ  �       �                    �?���}D�?-            �P@ �aQ  �       �                    �? ��WV�?             :@ 7aQ  ������������������������       �                     @       �       �                    6@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@       �       �                    @��]�T��?            �D@�aQ  �       �                    �?\�Uo��?             C@ saQ  ������������������������       �                      @EaQ  �       �                    @�q�q�?             B@�aQ  �       �                 03{3@�q�����?             9@        �       �                     @z�G�z�?             $@ aQ  �       �                    *@z�G�z�?             @ �aQ  ������������������������       �                     �?�aQ  ������������������������       �                     @ �aQ  �       �                   �5@z�G�z�?             @�aQ  ������������������������       �                     @iaQ  ������������������������       �                     �?        �       �                 �̌4@�q�q�?             .@ �aQ  ������������������������       �                     @       �       �                    �?�q�q�?             (@eaQ  �       �                    :@�z�G��?             $@       �       �                     @      �?             @        ������������������������       �                      @        �       �                    +@      �?              @ 4aQ  ������������������������       �                     �?       ������������������������       �                     �?�aQ  ������������������������       �                     @       ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                     @ 6aQ  �       �                 pf�C@�q�q�?             @        �       �                    @�q�q�?             @        ������������������������       �                      @aQ  ������������������������       �                     �? eaQ  ������������������������       �                     @       ������������������������       �                     @       �       �                    �?ƆQ����?P            �^@�aQ  �       �                  "�b@pY���D�?0            �S@       ������������������������       �        %            �M@        �       �                    �?ףp=
�?             4@�aQ  ������������������������       �                     $@       �       �                    $@z�G�z�?             $@ aQ  ������������������������       �                      @�aQ  ������������������������       �                      @        �                           @�&!��?             �E@       �                          �?p�ݯ��?             C@paQ  �                           �?b�2�tk�?             B@       �       	                �UwR@���Q��?            �A@ �aQ  �                          �?�<ݚ�?             2@                                  �?���Q��?             @        ������������������������       �                      @                             ��UO@�q�q�?             @       ������������������������       �                      @       ������������������������       �                     �?                               �C@$�q-�?             *@        ������������������������       �                     @                                F@؇���X�?             @        ������������������������       �                     �?       ������������������������       �                     @       
                         �?j���� �?             1@                                 �?      �?              @� ��t�                          �?؇���X�?             @                                �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                                �?z�G�z�?             @                              �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @                                =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @              $                p�O@���Q��?             @              #                   >@      �?             @       !      "                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�b�[     h�h*h-K ��h/��R�(KM%KK��h]�BP       �z@     �q@     �x@      h@      O@      `@      �?      0@              &@      �?      @      �?                      @     �N@      \@      @     �O@      @      5@      �?      (@              (@      �?               @      "@      �?       @      �?       @      �?                       @              @      �?      �?      �?                      �?      �?      E@              ?@      �?      &@              @      �?      @      �?                      @     �L@     �H@       @      (@       @      @       @       @               @       @                      @              @     �K@     �B@      <@      ?@      :@      1@      @      @      @                      @      7@      $@              @      7@      @      .@      @      @              $@      @      @      �?       @      �?       @                      �?      @              @      @      �?               @      @              @       @               @               @      ,@      �?              �?      ,@      �?       @      �?                       @              (@      ;@      @      3@       @               @      3@               @      @              �?       @      @      @              @      @       @              @      @       @      @              @       @              �?             �t@     @P@      `@      @     @^@      @      W@      @      A@      @      .@              3@      @               @      3@      @      "@              $@      @              �?      $@       @       @       @       @              M@       @      3@             �C@       @     �C@      �?      5@              2@      �?              �?      2@                      �?      =@               @             �i@      M@      @@      0@      �?      @               @      �?      @              @      �?              ?@      $@      <@      $@      .@      $@      @      "@      @      @      @      @               @      @      �?              �?      @              @      �?      �?      �?              �?      �?               @                      @      "@      �?      "@                      �?      *@              @             �e@      E@     @]@      2@     �G@      @      �?              G@      @     �F@      @      ?@      @      $@              5@      @      *@               @      @      @      @              �?      @       @       @              �?       @      @              ,@              �?             �Q@      .@      @             �P@      .@      @      @      @               @      @               @       @      @      �?       @      �?      �?     �N@      $@              �?     �N@      "@      8@      @      @      @              @      @              3@      @      .@      @      *@       @      @       @       @              @       @      @                       @      @               @       @       @                       @      @             �B@       @      5@       @      ,@              @       @      @      �?              �?      @                      �?      0@              L@      8@      @       @      �?       @      �?      @               @      �?      �?      �?                      �?              @      @             �I@      0@      9@      �?      @              6@      �?              �?      6@              :@      .@      7@      .@       @              5@      .@      (@      *@       @       @      �?      @      �?                      @      �?      @              @      �?              $@      @      @              @      @      @      @      �?      @               @      �?      �?              �?      �?              @                       @      "@       @      @              @       @      �?       @               @      �?              @              @              <@     �W@       @     @S@             �M@       @      2@              $@       @       @       @                       @      :@      1@      8@      ,@      6@      ,@      5@      ,@      ,@      @       @      @               @       @      �?       @                      �?      (@      �?      @              @      �?              �?      @              @      $@       @      @      �?      @      �?       @      �?                       @              @      �?              @      @      @      �?      �?      �?      �?                      �?      @              �?      @      �?      �?              �?      �?                       @      �?               @               @      @      �?      @      �?      �?              �?      �?                       @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJQY%hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @��ϙLq�?�           8�@               	                    @     ��?             @@ l                                @��.k���?             1@�aQ                             �?ףp=
�?             $@ �aQ                               @      �?              @ �aQ  ������������������������       �                     �?�aQ  ������������������������       �                     �?"5bQ  ������������������������       �                      @�aQ  ������������������������       �                     @        
                           �?��S�ۿ?
             .@       ������������������������       �                     $@       @                           @z�G�z�?             @      @������������������������       �                     @                                   �?      �?              @      $@������������������������       �                     �?      "@������������������������       �                     �?       @       �                 `fK@�ĸۦ��?�           8�@     (@       Q                    �?��J��?r           @�@               "                     @Z�2�t��?h            �d@               !                    �?0)RH'�?(            @Q@     @                          �*@�q�q��?             H@     @P@                           B@���Q��?             4@     @                          �9@      �?	             0@      @                          �'@z�G�z�?             @       @������������������������       �                     �?        ������������������������       �                     @      �?������������������������       �                     &@        ������������������������       �                     @      @                        ���;@ �Cc}�?             <@       ������������������������       �                     6@      "@                         X��C@      �?             @     �?������������������������       �                     @      �?������������������������       �                     @       @������������������������       �                     5@      �?#       0                 pF @�W*��?@            @X@        $       /                    �?��hJ,�?             A@       %       .                 X��B@<���D�?            �@@     4@&       '                   �6@     ��?             @@      $@������������������������       �                     .@        (       )                   �8@@�0�!��?             1@      3@������������������������       �                      @      @*       -                 ���@��S�ۿ?             .@      �?+       ,                 �Y�@      �?             @      �?������������������������       �                     @       @������������������������       �                     �?        ������������������������       �        	             &@      @������������������������       �                     �?      @������������������������       �                     �?      �?1       N                 03�7@����X�?+            �O@       2       K                    �?�D����?             E@     "@3       F                    �?p�ݯ��?             C@       4       ?                 ��.@     ��?             @@      @5       >                    �?�J�4�?             9@     �?6       ;                 �&�%@������?             1@       7       :                 `��!@ףp=
�?             $@      �?8       9                 `�X!@      �?             @     @������������������������       �                     @      �?������������������������       �                     �?       @������������������������       �                     @      �?<       =                 ���*@և���X�?             @        ������������������������       �                     @      &@������������������������       �                     @        ������������������������       �                      @        @       A                    �?؇���X�?             @      �?������������������������       �                     @      �?B       C                 03�1@      �?             @      �?������������������������       �                      @      @D       E                    �?      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      @G       J                    @�q�q�?             @      @H       I                   �4@���Q��?             @      @������������������������       �                      @       @������������������������       �                     @        ������������������������       �                     �?        L       M                 �|Y=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        O       P                    �?���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        R       �                   �J@T�1!�}�?
            z@       S       \                   �2@      �?�            �x@        T       [                 �&@������?             B@        U       V                    �?�X�<ݺ?             2@       ������������������������       �                     $@        W       Z                    �?      �?              @        X       Y                  �K"@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ]       x                     �?4�<����?�            @v@        ^       e                 �|�<@��J�fj�?            �B@        _       `                    7@      �?              @        ������������������������       �                     �?        a       b                 `f�D@؇���X�?             @       ������������������������       �                     @        c       d                 ��I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       w                   �G@J�8���?             =@       g       r                 �TA@@l��
I��?             ;@       h       m                 ���=@j���� �?             1@       i       l                 ��";@"pc�
�?
             &@       j       k                 ��:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        n       o                  �>@r�q��?             @        ������������������������       �                     @        p       q                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �C@ףp=
�?             $@       ������������������������       �                     @        u       v                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                    �?0�\>��?�            �s@       z       �                   @E@�u����?�             q@       {       �                    �?Ǖi�7�?�            0p@       |       �                     @X�EQ]N�?�             p@        }       ~                    �?���c���?             J@        ������������������������       �                     @               �                   @D@؇���X�?            �H@       �       �                 `fF)@�����H�?            �F@        �       �                    5@���7�?             6@ 910,15.������������������������       �                     �? 58,,S
6������������������������       �                     5@ 0.5,,S
�       �                 �|�<@�㙢�c�?             7@ rgue)",������������������������       �                      @ iss. El�       �                   �3@������?             .@,"Ander�       �                   �A@�	j*D�?             *@ale,39,�       �                    @@      �?              @,,0,0,S�       �                 �|�=@      �?             @  Jane",������������������������       �                     �? e,,0,0,������������������������       �                     @ male,35������������������������       �      �?             @ 24,1,2,������������������������       �                     @ 1,1,347������������������������       �                      @K Stanl������������������������       �      �?             @ss. Mar�       �                 �Y�@�"�_*d�?�            �i@ r. Lawr�       �                   �8@���y4F�?             C@ oni",ma�       �                   �3@���|���?             &@ son Jr"������������������������       �                     @id",male�       �                    5@      �?              @ ard",ma�       �                    �?�q�q�?             @  ""Dai"������������������������       �                      @ick",mal������������������������       �                     �?les Leo������������������������       �                     @ Gretch�       �                 ���@ 7���B�?             ;@ndyeff,������������������������       �                     6@nnell, ������������������������       �z�G�z�?             @rth, Mr�       �                 �?�@4և����?k             e@,3,"Lun�       �                 �?$@x��B�R�?9            �V@ 3,1,1,"�       �                    ;@�8��8��?             B@ 34,0,1,������������������������       �                     *@ ,0,3,"S�       �                  s�@�LQ�1	�?             7@ avis, M������������������������       �                     @ Mr. Ant�       �                    �?     ��?             0@,"Colly�       �                 �|Y=@"pc�
�?	             &@ Panula,������������������������       �                     �? .6875,,�       �                 X��A@ףp=
�?             $@6.1,,S
������������������������       ������H�?             "@ 2,,S
64������������������������       �                     �? B35,C
6�       �                 �|Y>@z�G�z�?             @ 8,27.9,������������������������       �      �?              @ 5,1,3,"������������������������       �                     @ 46,1,1,������������������������       �                    �K@ D33,C
6�       �                    �?� ���?2            @S@ 48,1,1,������������������������       �                     @35.5,A26�       �                   @C@�MI8d�?/            �R@.55,,S
�       �                   �3@؇���X�?,            �Q@ A. 2314������������������������       ����Q��?             @958,,S
�       �                 ��) @�?�<��?*            @P@653,0,3�       �                   �>@��(\���?             D@,,S
654������������������������       �                     =@,7.8292�       �                   �@@���!pc�?             &@0,36522�       �                   �?@      �?             @ ,S.O.C.������������������������       �                     �?349223,������������������������       ����Q��?             @32,1,1,������������������������       �                     @ e,23,0,�       �                 �|�>@z�G�z�?             9@8,0,2,3�       �                   �8@      �?             4@ ",male,������������������������       �                     @e,40,0,�       �                 0S%"@     ��?             0@ ,47,0,0�       �                 �|Y<@���Q��?             @ 0,34921������������������������       �                      @,1,0,ST�       �                 pf� @�q�q�?             @ e,32,2,������������������������       �                     �?on",mal������������������������       �                      @ ",male,�       �                   �<@"pc�
�?             &@ 0,A/5 3������������������������       �                     @ummins W�       �                 �|Y=@���Q��?             @ Thomas �       �                 ���"@�q�q�?             @ ,29750,������������������������       �                     �?2750,52������������������������       �                      @C.A. 24������������������������       �                      @ 44270,1������������������������       �                     @ 6,0,,S
�       �                   @D@      �?             @12,7.77�       �                 ��	0@�q�q�?             @ 0,34282������������������������       �                      @ ,4138,9������������������������       �                     �?",femal������������������������       �                     �? ke Mart������������������������       �                     �? ,"Peter������������������������       �                     .@ sab, Mr�       �                 ��.@`Ӹ����?            �F@ vigen, �       �                    �?r�q��?	             (@dwin, M�       �                     @�C��2(�?             &@ rown, M������������������������       �                     �? 2,"Laro�       �                    5@ףp=
�?             $@ 2123,41������������������������       �                     �?101295,������������������������       �                     "@,10.170������������������������       �                     �? 0,35003������������������������       �                    �@@ emale,1������������������������       �                     :@ n",male�       �                    �?�"�q��?A            �W@e,4,0,1�       �                    �?�}�+r��?'            �L@56.4958������������������������       �                     =@695,0,1�       �                    @ �Cc}�?             <@hapman,������������������������       �                     9@elly, M������������������������       �                     @ss. Kat�       �                    �?p�ݯ��?             C@ayer, M�       �                 X�,@@��Q��?             4@,"Humbl�       �                  �}S@      �?             $@ .65,F G������������������������       �                     @ Force)"�       �                    �?r�q��?             @thorne,������������������������       �                     @ 03,0,3,�       �                   �5@      �?              @ ,0,3,"G������������������������       �                     �?,"Hanse������������������������       �                     �?"Morley�       �                    �?z�G�z�?             $@50655,2�       �                   @H@�����H�?             "@0,0,223������������������������       �                     @male,42,�       �                   �T@�q�q�?             @ ,female������������������������       �                      @  Gonios������������������������       �                     �?,"Mayne,������������������������       �                     �?,0,PC 1�       �                     @b�2�tk�?             2@,113028�       �                     �?      �?	             (@1,0,199�       �                 �|Y>@�eP*L��?             &@ ,0,0,75������������������������       �                     �? 250647,�       �                    �?���Q��?             $@",male,�       �                 03�U@      �?              @e Louis�       �                    C@�q�q�?             @ Miss. E������������������������       �                     �?19,0,3,������������������������       �                      @hnson, ������������������������       �                     @,"Harper������������������������       �                      @722,0,3������������������������       �                     �?
723,0,�       �                    @r�q��?             @724,0,2������������������������       �                     @ ,1,"Cha������������������������       �                     �? 726,0,3�t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �|@     �o@      "@      7@       @      "@      �?      "@      �?      �?      �?                      �?               @      @              �?      ,@              $@      �?      @              @      �?      �?      �?                      �?     �{@      m@     �z@     @c@     �N@     @Z@      &@      M@      &@     �B@       @      (@      @      (@      @      �?              �?      @                      &@      @              @      9@              6@      @      @              @      @                      5@      I@     �G@      @      =@      @      =@      @      =@              .@      @      ,@       @              �?      ,@      �?      @              @      �?                      &@      �?              �?             �F@      2@      9@      1@      8@      ,@      6@      $@      5@      @      *@      @      "@      �?      @      �?      @                      �?      @              @      @              @      @               @              �?      @              @      �?      @               @      �?      �?      �?                      �?       @      @       @      @       @                      @              �?      �?      @              @      �?              4@      �?              �?      4@             w@     �H@     pu@     �H@     �A@      �?      1@      �?      $@              @      �?      @      �?      @                      �?      @              2@             @s@      H@      5@      0@       @      @      �?              �?      @              @      �?      �?      �?                      �?      3@      $@      3@       @      $@      @      "@       @      @       @      @                       @      @              �?      @              @      �?       @      �?                       @      "@      �?      @              @      �?      @                      �?               @     �q@      @@     �n@      >@     �l@      >@     �l@      >@     �F@      @      @              E@      @      D@      @      5@      �?              �?      5@              3@      @       @              &@      @      "@      @      @      @      @      �?              �?      @              �?      @      @               @               @       @     �f@      7@      >@       @      @      @      @              �?      @      �?       @               @      �?                      @      :@      �?      6@              @      �?      c@      .@      V@      @     �@@      @      *@              4@      @      @              *@      @      "@       @              �?      "@      �?       @      �?      �?              @      �?      �?      �?      @             �K@             @P@      (@      @              O@      (@      N@      $@      @       @     �L@       @     �B@      @      =@               @      @      @      @              �?      @       @      @              4@      @      .@      @      @              &@      @       @      @               @       @      �?              �?       @              "@       @      @              @       @      �?       @      �?                       @       @              @               @       @      �?       @               @      �?              �?              �?              .@             �E@       @      $@       @      $@      �?      �?              "@      �?              �?      "@                      �?     �@@              :@              1@     �S@      @      K@              =@      @      9@              9@      @              ,@      8@      @      *@      @      @              @      @      �?      @              �?      �?      �?                      �?       @       @      �?       @              @      �?       @               @      �?              �?              @      &@      @      @      @      @      �?              @      @       @      @       @      �?              �?       @                      @       @              �?              �?      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��fbhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM5huh*h-K ��h/��R�(KM5��h|�B@M         F                    �?�u����?�           8�@                                   �?sYi9��?O            `a@                                    @\#r��?"            �N@     @                          �H@��<b�ƥ?             G@�aQ  ������������������������       �                     E@      M@                           J@      �?             @      �?������������������������       �                     �?        ������������������������       �                     @      @	                           �?�q�q�?
             .@       
                           �?X�Cc�?	             ,@                                �&�)@և���X�?             @        ������������������������       �                     @       ������������������������       �                     @                               `�@1@����X�?             @                                 @      �?             @        ������������������������       �                      @       ������������������������       �                      @      @������������������������       �                     @      @������������������������       �                     �?      @       E                 �U�X@�θ�?-            �S@      @       D                  �	U@��R[s�?*            �Q@      @       C                    �?��ga�=�?(            �P@     @       <                 ��<J@�'�`d�?'            �P@     @       9                    �?&y�X���?#             M@      @       6                    �?r�����?             �J@      @       5                 p�i@@��k=.��?            �G@              2                   `A@�I�w�"�?             C@              1                 �|�=@"pc�
�?            �@@    @U@                             �?d}h���?             <@                                0C�<@      �?              @     �I@������������������������       �                     �?      &@������������������������       �                     �?        !       (                    ;@���B���?             :@      @"       '                 ���@�8��8��?             (@     @#       $                 ��y@؇���X�?             @      @������������������������       �                     �?      7@%       &                   �7@r�q��?             @      @������������������������       �                     �?      @������������������������       �                     @      .@������������������������       �                     @      @)       *                 �|Y=@����X�?	             ,@      �?������������������������       �                     �?      �?+       ,                     @�θ�?             *@      (@������������������������       �                     �?       @-       0                   @@      �?             (@     @.       /                 ���@      �?              @        ������������������������       �                     �?      @������������������������       �և���X�?             @      �?������������������������       �                     @       @������������������������       �                     @        3       4                      @���Q��?             @       @������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@      �?7       8                 �&�)@r�q��?             @      K@������������������������       �                     �?        ������������������������       �                     @      @:       ;                ��k/@z�G�z�?             @        ������������������������       �                     �?      @������������������������       �                     @        =       B                 ���Q@      �?              @       >       A                    �?      �?             @     �??       @                    F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?      �?������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     �?      @������������������������       �                     @      �?������������������������       �                      @      @G                          �?��s�ɝ�?t           ��@      @H       �                    �?>4և���?"            |@     @I       z                    �?������?�            �w@       @J       g                   �9@z�G�z�?2            �R@        K       `                   �6@�û��|�?             7@       L       _                 8#B2@������?             1@       M       N                   �1@���|���?
             &@        ������������������������       �                     �?        O       X                   �4@���Q��?	             $@       P       Q                    �?      �?             @        ������������������������       �                     �?        R       W                    3@���Q��?             @       S       T                 P��@      �?             @        ������������������������       �                     �?        U       V                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                     @      �?             @        ������������������������       �                     �?        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ]       ^                 pF�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        a       b                     @r�q��?             @        ������������������������       �                     �?        c       f                    8@z�G�z�?             @       d       e                 @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                      @       h       i                    �?ȵHPS!�?!             J@        ������������������������       �                     $@       j       w                     @؇���X�?             E@       k       n                 `f&'@ >�֕�?            �A@        l       m                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        o       p                     �?�g�y��?             ?@        ������������������������       �                     *@        q       r                   �B@�X�<ݺ?             2@       ������������������������       �                     "@        s       v                   �*@�����H�?             "@        t       u                    D@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        x       y                 �|�;@և���X�?             @        ������������������������       �                     @       ������������������������       �                     @       {       �                 ��$:@�Qb��?�            �r@       |       �                   @@@������?�            0p@       }       �                   �>@$�3c�s�?v            �g@       ~       �                 @3�@��I�� �?o            `f@              �                 �|Y=@��<D�m�?;            �X@        �       �                 ��@      �?             D@       �       �                  ��@z�G�z�?             9@       �       �                    �?�C��2(�?             6@ i6bQ  ������������������������       �                     �?�w6bQ  �       �                    7@�����?             5@76bQ  ������������������������       �                     (@        �       �                 ���@�<ݚ�?             "@        �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @ a6bQ  ������������������������       �                     @ 26bQ  ������������������������       �                     @        ������������������������       �                     .@@;6bQ  �       �                 �|�=@ _�@�Y�?             M@       �       �                     @@3����?             K@        ������������������������       �                     &@        �       �                 ��@ qP��B�?            �E@       ������������������������       �                     6@t6bQ  �       �                 �Y5@���N8�?
             5@        ������������������������       �z�G�z�?             @       ������������������������       �                     0@        ������������������������       �                     @�6bQ  �       �                   �3@�
��P�?4            @T@ �6bQ  �       �                   �2@�d�����?             3@       �       �                 ��Y @ףp=
�?             $@ L6bQ  �       �                    1@      �?              @        ������������������������       �                     �?�<6bQ  ������������������������       �                     �?        ������������������������       �                      @�3bQ  �       �                 ���$@X�<ݚ�?             "@       �       �                 0S5 @����X�?             @        ������������������������       ��q�q�?             @ �6bQ  ������������������������       �                     @        ������������������������       �                      @       �       �                    �?��a�n`�?(             O@ �4bQ  ������������������������       �                     �?       �       �                 ��) @\#r��?'            �N@        ������������������������       �                     6@        �       �                    :@8�Z$���?            �C@ �3bQ  ������������������������       �                     .@        �       �                     @      �?             8@        �       �                 �|Y<@�8��8��?             (@        ������������������������       �                     @ �6bQ  �       �                     �?؇���X�?             @        ������������������������       �                      @�4bQ  �       �                 �|�=@z�G�z�?             @        ������������������������       �                     �?�U6bQ  ������������������������       �                     @ �6bQ  �       �                 0S%"@�q�q�?             (@        �       �                 pf� @z�G�z�?             @        ������������������������       �                      @�6bQ  �       �                 �|Y<@�q�q�?             @ �6bQ  ������������������������       �                      @ �4bQ  ������������������������       �                     �?        �       �                 �|�=@؇���X�?             @n6bQ  ������������������������       �                     @        ������������������������       �                     �?��6bQ  �       �                 �&B@X�<ݚ�?             "@        ������������������������       �                     �? �3bQ  �       �                   �@      �?              @ �3bQ  ������������������������       �                     @        �       �                 �?�@���Q��?             @ U6bQ  ������������������������       �                     �?`e6bQ  �       �                 ��I @      �?             @6bQ  �       �                   �?@�q�q�?             @ �4bQ  ������������������������       �                     �?       ������������������������       �      �?              @        ������������������������       �                     �?�=/bQ  �       �                   @E@�J�T�?-            �Q@6bQ  �       �                 �?�@�X�<ݺ?             B@        ������������������������       �        
             1@       �       �                 @3�@�KM�]�?             3@ S1bQ  ������������������������       ��q�q�?             @��6bQ  �       �                   @D@      �?             0@d6bQ  ������������������������       �                     ,@        �       �                     @      �?              @ 16bQ  ������������������������       �                     �?        ������������������������       �                     �?Pz6bQ  ������������������������       �                    �A@ 86bQ  �       �                     �?X��ʑ��?            �E@}6bQ  �       �                 ��yC@j���� �?             A@       �       �                   �A@����X�?             <@       �       �                 �T!@@�q�q�?             8@       �       �                   �J@���!pc�?             6@       �       �                 `fF<@�t����?	             1@,6bQ  �       �                 �|�?@$�q-�?             *@ 5bQ  ������������������������       �                     �?05bQ  ������������������������       �                     (@ �3bQ  �       �                   @>@      �?             @        ������������������������       �                     �?``6bQ  ������������������������       �                     @�4bQ  �       �                 `fF<@z�G�z�?             @6bQ  ������������������������       �                     @ +6bQ  ������������������������       �                     �?�W3bQ  ������������������������       �                      @0�3bQ  ������������������������       �                     @        ������������������������       �                     @P&6bQ  �       �                    ;@�<ݚ�?             "@        �       �                 ��?P@�q�q�?             @ �6bQ  ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     @       �       �                   �:@DX�\��?3            �Q@ z6bQ  �       �                    �?��2(&�?             6@       �       �                     @     ��?             0@ '6bQ  �       �                    2@����X�?             @        ������������������������       �                     �?        �       �                     �?r�q��?             @        ������������������������       �                      @�|6bQ  �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @ �3bQ  �       �                   �!@�����H�?             "@ �3bQ  �       �                 ��Y@      �?             @        ������������������������       �                     @       ������������������������       �                     �?�7bQ  ������������������������       �                     @        ������������������������       �                     @        �       �                    �?Rg��J��?%            �H@ C6bQ  �       �                   @C@���|���?             &@       �       �                    �?�z�G��?             $@T6bQ  ������������������������       �                     @ !6bQ  ������������������������       �                     @        ������������������������       �                     �?        �                           @      �?             C@�6bQ  �                         @D@��}*_��?             ;@       �                           �?�<ݚ�?             2@6bQ  �                       �|Y=@r�q��?	             (@                               ���M@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?                                �?ףp=
�?             $@       ������������������������       �                     @                              `f�K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �@@�q�q�?             @       	      
                  �<@z�G�z�?             @        ������������������������       �                     �?                                �7@      �?             @ � �q� ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �?�q�q�?             "@                             �CdQ@      �?              @        ������������������������       �                     @                                 �?���Q��?             @        ������������������������       �                      @                              ��#[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?"pc�
�?             &@                              ���.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              (                    @�^�����?R             _@                                 �? i���t�?$            �H@       ������������������������       �                     C@               !                   �?�eP*L��?             &@        ������������������������       �                     �?        "      '                   �?���Q��?             $@       #      $                    �?X�<ݚ�?             "@        ������������������������       �                      @        %      &                   :@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        )      4                   �?��n�?.            �R@        *      +                  �7@���Q��?            �A@        ������������������������       �                     (@        ,      1                ��T?@���}<S�?             7@       -      0                   @@�}�+r��?             3@        .      /                �|Y>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        2      3                ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@        �t�bh�h*h-K ��h/��R�(KM5KK��h]�BP       �{@     �p@     �P@     @R@      @     �K@      �?     �F@              E@      �?      @      �?                      @      @      $@      @      "@      @      @              @      @               @      @       @       @               @       @                      @              �?      N@      2@      J@      2@      J@      .@      J@      ,@     �G@      &@     �E@      $@      C@      "@      =@      "@      ;@      @      6@      @      �?      �?      �?                      �?      5@      @      &@      �?      @      �?      �?              @      �?              �?      @              @              $@      @              �?      $@      @      �?              "@      @      @      @      �?              @      @      @              @               @      @              @       @              "@              @      �?              �?      @              @      �?              �?      @              @      @      �?      @      �?      �?              �?      �?                       @      @                      �?              @       @             �w@      h@     �s@     �`@     �p@     �Z@      .@      N@      "@      ,@      @      *@      @      @              �?      @      @      @      @              �?      @       @       @       @              �?       @      �?       @                      �?      �?              �?      @              �?      �?       @              �?      �?      �?              �?      �?                      @      @      �?      �?              @      �?       @      �?              �?       @               @              @      G@              $@      @      B@       @     �@@      �?      @              @      �?              �?      >@              *@      �?      1@              "@      �?       @      �?      @      �?                      @              @      @      @              @      @              p@      G@     `m@      8@     �d@      6@     @d@      1@      W@      @     �A@      @      4@      @      4@       @      �?              3@       @      (@              @       @      �?       @      �?                       @      @                      @      .@             �L@      �?     �J@      �?      &@              E@      �?      6@              4@      �?      @      �?      0@              @             �Q@      &@      ,@      @      "@      �?      �?      �?      �?                      �?       @              @      @      @       @      �?       @      @                       @      L@      @      �?             �K@      @      6@             �@@      @      .@              2@      @      &@      �?      @              @      �?       @              @      �?              �?      @              @      @      �?      @               @      �?       @               @      �?              @      �?      @                      �?      @      @      �?              @      @              @      @       @      �?               @       @      �?       @              �?      �?      �?      �?             @Q@       @      A@       @      1@              1@       @       @      �?      .@      �?      ,@              �?      �?              �?      �?             �A@              5@      6@      ,@      4@       @      4@       @      0@      @      0@       @      .@      �?      (@      �?                      (@      �?      @      �?                      @      @      �?      @                      �?       @                      @      @              @       @      �?       @               @      �?              @              E@      =@      3@      @      *@      @      @       @              �?      @      �?       @              @      �?              �?      @               @      �?      @      �?      @                      �?      @              @              7@      :@      @      @      @      @              @      @              �?              3@      3@      $@      1@      @      ,@       @      $@      �?      �?              �?      �?              �?      "@              @      �?       @      �?                       @       @      @      �?      @              �?      �?      @      �?                      @      �?              @      @      @      @      @               @      @               @       @      �?       @                      �?      �?              "@       @      �?       @      �?                       @       @             �P@      M@      @      F@              C@      @      @      �?              @      @      @      @       @               @      @              @       @                      �?     �N@      ,@      5@      ,@              (@      5@       @      2@      �?      @      �?      @                      �?      ,@              @      �?              �?      @              D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ$�phG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         .                   �3@�L*�<�?�           8�@ d4bQ         +                    @b�L�4��?P            �`@     �?                           �?�Sb(�	�?A             [@       @                           �?���.�6�?             G@      @������������������������       �        
             2@     @                            @ �Cc}�?             <@     @������������������������       �                     2@      "@       	                    @�z�G��?             $@      �?������������������������       �                     @        
                           �?      �?             @                                  �?      �?             @       ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                      @                               �?�@�g�y��?#             O@        ������������������������       �                     ,@                                   �?      �?             H@      @������������������������       �                      @      @                            �?�LQ�1	�?             G@      @                           �?և���X�?             <@      @                            @      �?
             8@       @                          �2@      �?             @      @������������������������       �                      @     @                          �'@      �?             @       @������������������������       �                     @      @������������������������       �                     �?                               ��Y @      �?             2@                                  1@ףp=
�?             $@     @U@������������������������       �      �?             @        ������������������������       �                     @     �I@������������������������       �                      @      &@������������������������       �                     @        !       "                    �?�<ݚ�?             2@       @������������������������       �                      @        #       $                 03{3@      �?             0@        ������������������������       �                     $@      �?%       *                    �?�q�q�?             @       &       )                    �?���Q��?             @     �?'       (                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @      @������������������������       �                     �?      @������������������������       �                     �?        ,       -                   -@$�q-�?             :@      @������������������������       �                      @       @������������������������       �                     8@      �?/       p                    �?B�����?_           �@      @0       A                     @tHN�?q             f@      @1       >                   @L@X'"7��?H             [@      @2       3                    �?T��,��?D            @Y@      �?������������������������       �                     A@      �?4       =                    �?�����?-            �P@     4@5       6                   �B@@4և���?             E@     .@������������������������       �                     =@      @7       8                   @C@�θ�?	             *@        ������������������������       �                     �?        9       :                     �?r�q��?             (@        ������������������������       �                     @      @;       <                    �?����X�?             @       ������������������������       �                     @      �?������������������������       �                      @        ������������������������       �                     9@      @?       @                   �L@����X�?             @      3@������������������������       �                      @      �?������������������������       �                     @      @B       m                    @\X��t�?)            @Q@     @C       l                 03�:@p�EG/��?%            �O@       D       S                    �?d��0u��?"             N@      @E       R                    �?������?             >@     �?F       Q                 ��.@l��
I��?             ;@      @G       H                 �|Y=@X�<ݚ�?	             2@        ������������������������       �                     �?      @I       N                    �?��.k���?             1@        J       M                    �?�<ݚ�?             "@     �?K       L                 X�x&@�q�q�?             @       @������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     @        O       P                 �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        T       k                   @B@��S���?             >@       U       f                    �?�5��?             ;@       V       ]                    �?      �?             4@       W       Z                 ��� @��
ц��?             *@       X       Y                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                 ���)@և���X�?             @        ������������������������       �                      @        `       e                 03�1@���Q��?             @       a       d                   �0@      �?             @       b       c                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        g       h                    �?؇���X�?             @        ������������������������       �                     @        i       j                 �|�:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       o                 ���4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        q       �                 ��D:@\���(\�?�             y@       r       �                    �?\2R}�?�            r@        s       ~                 �|Y=@�θV�?,            @Q@        t       }                    �?����X�?
             ,@       u       z                    �?�q�q�?             (@       v       w                   �8@�z�G��?             $@        ������������������������       �                     @        x       y                   @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        {       |                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               �                 �|�=@�1�`jg�?"            �K@       �       �                    �?Du9iH��?            �E@        �       �                    �?$�q-�?
             *@910,15.������������������������       �        	             (@ 58,,S
6������������������������       �                     �? 0.5,,S
�       �                   `3@��S�ۿ?             >@rgue)",�       �                 ���@h�����?             <@ iss. El������������������������       �                     $@,"Ander�       �                   @'@�X�<ݺ?
             2@ale,39,������������������������       �$�q-�?             *@,,0,0,S������������������������       �                     @  Jane",�       �                    �?      �?              @ e,,0,0,������������������������       �                     �? male,35������������������������       �                     �? 24,1,2,������������������������       �                     (@ 1,1,347�       �                   @4@�2�~w�?�            �k@ K Stanl�       �                 pf� @      �?             0@ ss. Mar�       �                    �?      �?              @r. Lawr������������������������       �                     @ oni",ma������������������������       �                     @ son Jr"������������������������       �                      @id",male�       �                   �<@ =[y��?y            �i@ ard",ma������������������������       �        '            @P@  ""Dai"�       �                   �*@��X�-�?R            `a@ck",mal�       �                     @�#-���?@            @Z@ les Leo�       �                   �F@r�q��?             8@ Gretch�       �                   @D@���y4F�?             3@ndyeff,�       �                 `fF)@r�q��?             2@nnell, ������������������������       �                     $@rth, Mr�       �                 �|�=@      �?              @ ,3,"Lun������������������������       �                      @ 3,1,1,"�       �                    @@r�q��?             @ 34,0,1,������������������������       �                     @ ,0,3,"S�       �                   @B@�q�q�?             @avis, M������������������������       �      �?              @ Mr. Ant������������������������       �                     �?,"Colly������������������������       �                     �? Panula,������������������������       �                     @ .6875,,�       �                 ���"@xdQ�m��?/            @T@6.1,,S
�       �                 ��@ �\���?-            �S@ 2,,S
64������������������������       �                     7@ B35,C
6�       �                 ��L@@4և���?!             L@ 8,27.9,�       �                 �|Y>@���Q��?             @ 5,1,3,"������������������������       �                      @ 46,1,1,������������������������       �                     @ D33,C
6�       �                   �@@`'�J�?            �I@48,1,1,�       �                 ��) @`Jj��?             ?@5.5,A26�       �                 @3�@h�����?             <@.55,,S
�       �                 �?�@��S�ۿ?             .@A. 2314������������������������       �                     $@958,,S
������������������������       �z�G�z�?             @653,0,3������������������������       �                     *@,,S
654�       �                 �|Y=@�q�q�?             @ ,7.8292������������������������       �                     �?0,36522�       �                 �|�>@      �?              @ ,S.O.C.������������������������       �                     �?349223,������������������������       �                     �?32,1,1,������������������������       �        	             4@ e,23,0,�       �                    ?@      �?              @ 8,0,2,3������������������������       �                     �? ",male,������������������������       �                     �?e,40,0,������������������������       �                     A@ ,47,0,0�       �                 p�w@�/e�U��?A            �[@0,34921�       �                    �?� �W�??            �Z@,1,0,ST�       �                    �?X�Cc�?4             U@ e,32,2,�       �                 @�pX@
;&����?             7@on",mal�       �                    �?b�2�tk�?             2@",male,�       �                 �|�;@�eP*L��?             &@ 0,A/5 3������������������������       �                      @ummins W�       �                 ��2>@�q�q�?             "@ Thomas ������������������������       �                      @ ,29750,�       �                    C@؇���X�?             @2750,52������������������������       �                     @C.A. 24�       �                 �D D@�q�q�?             @ 44270,1������������������������       �                     �? 6,0,,S
������������������������       �                      @12,7.77�       �                 ��`E@؇���X�?             @ 0,34282������������������������       �                     �? ,4138,9������������������������       �                     @",femal������������������������       �                     @ ke Mart�       �                    R@�ɞ`s�?%            �N@,"Peter�       �                 03k:@�c�Α�?$             M@ sab, Mr������������������������       �                      @ vigen, �       �                 �!fK@      �?#             L@dwin, M�       �                     �?z�G�z�?             D@rown, M�       �                    <@��G���?            �B@ 2,"Laro������������������������       �                     �? 2123,41�       �                   �F@r�q��?             B@101295,�       �                    �?�E��ӭ�?             2@,10.170�       �                   `@@�n_Y�K�?
             *@ 0,35003�       �                 �|Y=@r�q��?             @ emale,1������������������������       �                     �? n",male������������������������       �                     @e,4,0,1������������������������       �                     @56.4958������������������������       �                     @695,0,1�       �                   @J@�X�<ݺ?
             2@ hapman,�       �                 `f�;@      �?              @ elly, M������������������������       �                     �?ss. Kat������������������������       �                     @ayer, M������������������������       �                     $@,"Humbl������������������������       �                     @ .65,F G�       �                    �?     ��?             0@Force)"�       �                     @�n_Y�K�?	             *@thorne,�       �                    C@�<ݚ�?             "@03,0,3,�       �                 �|Y>@���Q��?             @,0,3,"G������������������������       �                     @,"Hanse������������������������       �                      @"Morley������������������������       �                     @50655,2�       �                    >@      �?             @0,0,223�       �                    ;@      �?              @ ale,42,������������������������       �                     �? ,female������������������������       �                     �?  Gonios������������������������       �                      @,"Mayne,�       �                 ���[@�q�q�?             @ ,0,PC 1������������������������       �                     �?,113028������������������������       �                      @1,0,199������������������������       �                     @ ,0,0,75�       �                     �?�nkK�?             7@250647,�       �                    �?�8��8��?             (@ ",male,�       �                 ��UO@؇���X�?             @ e Louis������������������������       �                     @ Miss. E�       �                   @D@�q�q�?             @ 19,0,3,������������������������       �                     �?hnson, ������������������������       �                      @,"Harper������������������������       �                     @722,0,3������������������������       �                     &@
723,0,������������������������       �                     @724,0,2�t�b�     h�h*h-K ��h/��R�(KK�KK��h]�B�       p{@      q@     �M@     �R@     �A@     @R@      @     �E@              2@      @      9@              2@      @      @              @      @      @      �?      @              @      �?               @              @@      >@      ,@              2@      >@       @              0@      >@      (@      0@      (@      (@      @      @       @              �?      @              @      �?              "@      "@      �?      "@      �?      @              @       @                      @      @      ,@       @               @      ,@              $@       @      @       @      @       @       @       @                       @              �?              �?      8@       @               @      8@             �w@     �h@     �A@     �a@      @     �Y@      @     �X@              A@      @      P@      @     �C@              =@      @      $@      �?               @      $@              @       @      @              @       @                      9@       @      @       @                      @      >@     �C@      9@      C@      6@      C@       @      6@       @      3@       @      $@              �?       @      "@      @       @      @       @               @      @              @              �?      @      �?                      @              "@              @      ,@      0@      &@      0@      $@      $@      @      @      @       @               @      @              �?      @      �?                      @      @      @       @               @      @      �?      @      �?      �?      �?                      �?               @      �?              �?      @              @      �?       @               @      �?              @              @              @      �?              �?      @             �u@     �K@     �p@      4@      O@      @      $@      @       @      @      @      @      @              �?      @      �?                      @      �?      �?      �?                      �?       @              J@      @      D@      @      (@      �?      (@                      �?      <@       @      ;@      �?      $@              1@      �?      (@      �?      @              �?      �?      �?                      �?      (@             �i@      *@      (@      @      @      @      @                      @       @             `h@      "@     @P@             @`@      "@      X@      "@      4@      @      .@      @      .@      @      $@              @      @               @      @      �?      @               @      �?      �?      �?      �?                      �?      @              S@      @     �R@      @      7@              J@      @      @       @               @      @             �H@       @      =@       @      ;@      �?      ,@      �?      $@              @      �?      *@               @      �?      �?              �?      �?              �?      �?              4@              �?      �?              �?      �?              A@              S@     �A@      S@      ?@      K@      >@      (@      &@      @      &@      @      @               @      @      @               @      @      �?      @               @      �?              �?       @              �?      @      �?                      @      @              E@      3@      E@      0@               @      E@      ,@     �@@      @      >@      @              �?      >@      @      *@      @       @      @      �?      @      �?                      @      @              @              1@      �?      @      �?              �?      @              $@              @              "@      @       @      @      @       @      @       @      @                       @      @              �?      @      �?      �?              �?      �?                       @      �?       @      �?                       @              @      6@      �?      &@      �?      @      �?      @               @      �?              �?       @              @              &@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW:+LhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         r                    �?]@f�
�?�           8�@               a                    �?��K�"�?�            �q@      @       &                 `f�$@�e�U��?�            �m@       @       %                    �?��H�}�?              I@     @       "                    �?(���@��?            �G@     2@                        �̌@���� �?            �D@     &@                        ���@�r����?             >@      @       	                 �|Y:@����X�?             @      �?������������������������       �                     @        
                           �?�q�q�?             @ ���n	 �������������������������       �                     �?        ������������������������       �                      @  �?  �?                           �?���}<S�?             7@3�@33�@������������������������       �        	             0@��
AffA                           4@����X�?             @  HB  `B������������������������       �                     �?                                �&B@r�q��?             @     C@                          �7@�q�q�?             @      �?������������������������       �                      @       @������������������������       �                     �?        ������������������������       �                     @      0@                          �2@���|���?             &@       @������������������������       �                     �?                                ��� @�z�G��?             $@     @                        @3�@r�q��?             @     �?                          �8@�q�q�?             @      @������������������������       �                     �?                                   ;@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      @������������������������       �                     @                !                  SE"@      �?             @      @������������������������       �                      @      0@������������������������       �                      @      "@#       $                   �3@�q�q�?             @      @������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     @      0@'       `                 �QD@X�E)9�?v            �g@     *@(       E                    �?�<�}���?K            @^@     @)       D                    @�? Da�?(            �O@      @*       +                    �?\#r��?&            �N@        ������������������������       �                     @      @,       5                 `f�)@ �Cc}�?#             L@      �?-       .                 pF%@`2U0*��?             9@      @������������������������       �                     *@      �?/       0                    +@�8��8��?             (@      @������������������������       �                     @      �?1       4                    �?r�q��?             @      @2       3                 ��&@z�G�z�?             @      �?������������������������       �                     �?      �?������������������������       �                     @      �?������������������������       �                     �?      �?6       =                   �*@�חF�P�?             ?@      �?7       <                   �B@X�<ݚ�?             "@     4@8       ;                    �?����X�?             @     (@9       :                    <@�q�q�?             @      @������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     �?      @������������������������       �                      @      �?>       ?                    �?���7�?             6@     @������������������������       �                     .@        @       C                    1@؇���X�?             @       A       B                    "@�q�q�?             @     @������������������������       �                      @     @������������������������       �                     �?       ������������������������       �                     @      @������������������������       �                      @     �?F       _                   �@@V�a�� �?#             M@      @G       H                    �?F�t�K��?"            �L@        ������������������������       �        	             .@      @I       J                   �9@0,Tg��?             E@        ������������������������       �                     ,@     �?K       T                     @��>4և�?             <@      @L       M                    6@      �?             0@      �?������������������������       �                      @        N       S                    :@؇���X�?
             ,@       O       P                   �8@�<ݚ�?             "@        ������������������������       �                     �?        Q       R                   �E@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @       U       ^                 �̤=@�q�q�?             (@       V       ]                 `fV6@�z�G��?             $@       W       X                 �|�;@և���X�?             @        ������������������������       �                     @        Y       Z                 03�1@      �?             @        ������������������������       �                      @        [       \                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �        +             Q@       b       q                    @v�2t5�?            �D@       c       d                    �?      �?             A@        ������������������������       �                     @        e       f                     @�f7�z�?             =@        ������������������������       �                     @        g       h                    @�q�q�?             8@        ������������������������       �                     @        i       n                    *@p�ݯ��?
             3@       j       k                    @�8��8��?             (@        ������������������������       �                     @        l       m                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        o       p                 ���4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                     @        s       �                 ��D:@���<��?           �z@       t       y                    $@�%�P��?�            �t@        u       v                     @"pc�
�?             &@        ������������������������       �                     @        w       x                 ��|2@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        z       �                     @ E�+0+�?�            �s@        {       |                   �)@�(\����?1             T@        ������������������������       �                    �A@        }       �                 ��,@`Ӹ����?            �F@       ~                        �|�<@$�q-�?             :@        ������������������������       �                     ,@       �       �                 �|�=@r�q��?             (@        ������������������������       �                     �?        �       �                   �A@�C��2(�?             &@       �       �                    @@r�q��?             @        ������������������������       �                      @       ������������������������       �      �?             @        ������������������������       �                     @       ������������������������       �                     3@        �       �                    �?��5Վ3�?�            �m@        �       �                    �?^������?            �A@       �       �                    �?�c�Α�?             =@       �       �                 ���@      �?             8@        ������������������������       �                     @        �       �                   @@�q�q�?
             2@        �       �                   �5@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �|=@և���X�?             @        ������������������������       �                      @       ������������������������       ����Q��?             @        �       �                 �|�;@�����H�?             "@        �       �                   �2@      �?             @        ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                     @        �       �                 �&�)@���Q��?             @        ������������������������       �                      @       ������������������������       �                     @        �       �                 ��y&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@@ ��fί�?�            `i@       �       �                    �?3��e��?j            �d@       �       �                   �:@$s��O�?Z            �a@        �       �                   �2@�FVQ&�?,            �P@        �       �                   �1@      �?
             (@       �       �                   �0@�<ݚ�?             "@       �       �                 pf�@����X�?             @        ������������������������       �                      @       �       �                 pFD!@���Q��?             @        ������������������������       ��q�q�?             @       ������������������������       �                      @       ������������������������       �                      @        �       �                 ���@�q�q�?             @        ������������������������       �                     �?       �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@3����?"             K@        ������������������������       �                      @        �       �                 ���@ pƵHP�?!             J@        �       �                    7@z�G�z�?             @        ������������������������       �                      @        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                    �G@        �       �                 ��) @��A��?.            �R@       �       �                 @3�@lGts��?$            �K@       �       �                   �>@(L���?            �E@       �       �                 �|Y=@     ��?             @@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��(@�>����?             ;@       �       �                 03�@      �?             0@        ������������������������       �                     @       ������������������������       �"pc�
�?             &@        ������������������������       �                     &@       �       �                   �?@���!pc�?             &@        �       �                 pff@�q�q�?             @        ������������������������       �                     @       ������������������������       �                      @        �       �                 �?�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     (@        �       �                 ��)"@p�ݯ��?
             3@        �       �                 �|Y<@      �?              @        ������������������������       �                     @        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        �       �                    �?�C��2(�?             &@        ������������������������       �                      @       �       �                    (@�����H�?             "@        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        ������������������������       �                     @       �       �                    �? 7���B�?             ;@       ������������������������       �                     6@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     B@        �                          �J@*Mp����?J            �Y@       �       �                 ��";@|jq��?<            �T@        �       �                 03k:@      �?              @        ������������������������       �                     �?        �       �                 �|�?@����X�?             @        ������������������������       �                     �?       �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                   �C@      �?             @        ������������������������       �                     �?       �       �                    H@�q�q�?             @       ������������������������       �      �?              @       ������������������������       �                     �?        �       �                   �;@L�qA��?5            �R@        �       �                    6@l��[B��?             =@       �       �                    �?�����?             3@       ������������������������       �                     "@       �       �                    @���Q��?             $@        ������������������������       �                     @        �       �                    @�q�q�?             @       �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �                           �?���j��?!             G@       �                         �I@P����?             C@       �                          �?<ݚ)�?             B@       �                         �H@����X�?            �A@                              p�w@     ��?             @@                                �?������?             >@                             `f�B@�GN�z�?             6@                               �A@�eP*L��?	             &@             	                   �?�q�q�?             "@                              �|�=@�q�q�?             @        ������������������������       �                     �?                                �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       
                        �>@r�q��?             @                               @=@�q�q�?             @ � +�q� ������������������������       �                     �?                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                                 �?      �?              @                             `ށK@և���X�?             @        ������������������������       �                      @                                �G@���Q��?             @                                @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        !      (                   �?�}�+r��?             3@       "      #                   �?$�q-�?	             *@        ������������������������       �                     @        $      '                 )?@r�q��?             @        %      &                  �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       z@     `r@      O@     @k@      C@      i@      2@      @@      .@      @@      &@      >@      @      :@       @      @              @       @      �?              �?       @               @      5@              0@       @      @      �?              �?      @      �?       @               @      �?                      @      @      @              �?      @      @      @      �?       @      �?      �?              �?      �?              �?      �?              @               @       @               @       @              @       @               @      @              @              4@      e@      4@     @Y@       @     �K@      @     �K@              @      @      I@      �?      8@              *@      �?      &@              @      �?      @      �?      @      �?                      @              �?      @      :@      @      @       @      @       @      @       @                      @              �?       @              �?      5@              .@      �?      @      �?       @               @      �?                      @       @              (@      G@      &@      G@              .@      &@      ?@              ,@      &@      1@      @      (@       @               @      (@       @      @              �?       @      @              @       @                      @      @      @      @      @      @      @      @              �?      @               @      �?      �?      �?                      �?      @                       @      �?                      Q@      8@      1@      1@      1@              @      1@      (@              @      1@      @      @              (@      @      &@      �?      @              @      �?              �?      @              �?      @              @      �?              @             0v@      S@      r@     �D@       @      "@              @       @      @              @       @             �q@      @@     �S@       @     �A@             �E@       @      8@       @      ,@              $@       @              �?      $@      �?      @      �?       @              @      �?      @              3@              j@      >@      7@      (@      5@       @      2@      @      @              (@      @      @      @               @      @      @       @               @      @       @      �?      @      �?      @                      �?      @              @       @               @      @               @      @       @                      @      g@      2@     �b@      2@     �^@      1@      O@      @      "@      @      @       @      @       @       @              @       @      �?       @       @               @               @      �?      �?              �?      �?              �?      �?             �J@      �?       @             �I@      �?      @      �?       @               @      �?              �?       @             �G@             �N@      *@     �H@      @     �B@      @      =@      @      @      �?              �?      @              9@       @      ,@       @      @              "@       @      &@               @      @      @       @      @                       @      @      �?       @               @      �?      (@              (@      @       @      @              @       @      �?              �?       @              $@      �?       @               @      �?      @      �?       @               @      �?              �?       @              @              :@      �?      6@              @      �?              �?      @              B@             �P@     �A@     �H@      A@       @      @              �?       @      @      �?              �?      @               @      �?      @              �?      �?       @      �?      �?              �?     �G@      <@      ,@      .@      *@      @      "@              @      @              @      @       @      @       @               @      @              �?              �?      "@              "@      �?             �@@      *@      9@      *@      9@      &@      9@      $@      6@      $@      6@       @      1@      @      @      @      @      @      �?       @              �?      �?      �?      �?                      �?      @      �?       @      �?      �?              �?      �?      �?                      �?      @                       @      &@              @      @      @      @       @               @      @       @      �?              �?       @                       @      �?                       @      @                      �?               @       @              2@      �?      (@      �?      @              @      �?      �?      �?      �?                      �?      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJF<KdhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM'huh*h-K ��h/��R�(KM'��h|�B�I                             @	dm#��?�           8�@                                   @     ��?              H@     A@                        �-]@(;L]n�?             >@      @������������������������       �                     <@     @                        �(\�?      �?              @      M@������������������������       �                     �?      �?������������������������       �                     �?               	                    �?�<ݚ�?
             2@      @������������������������       �                     $@      @
                        ��T?@      �?              @      �?������������������������       �                      @      �?                           @�q�q�?             @     �?������������������������       �                     @      �?������������������������       �                      @       @       "                  @L@^ɼ���?�           ��@      @       W                    �?@\L5�T�?�           ؃@       @       4                     @l��TO��?H            @_@     C@                           �?�M���?(             Q@      �?                        03�=@�X�<ݺ?             B@       @                            �?      �?              @        ������������������������       �                      @      0@������������������������       �                     @       @������������������������       �                     <@               )                 �D�G@     ��?             @@     @                          �;@��.k���?             1@      �?������������������������       �                     �?      @       (                     �?     ��?
             0@              '                    �?��
ц��?             *@              &                    C@�q�q�?             (@     @       %                   �A@�eP*L��?             &@     @       $                 ��2>@���Q��?             $@               #                 �ܵ<@      �?              @     @!       "                 X�,@@      �?             @      @������������������������       �                      @       @������������������������       �                      @       @������������������������       �                     @      $@������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                     �?      @������������������������       �                     �?      :@������������������������       �                     @       @*       +                  �}S@������?
             .@      �?������������������������       �                     @      &@,       3                    �?      �?              @      @-       2                    �?�q�q�?             @      @.       1                    �?      �?             @     �?/       0                   �=@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @       @������������������������       �                     �?      �?������������������������       �                      @      @������������������������       �                      @      P@5       N                    �?�MWl��?             �L@     @6       9                    �?:	��ʵ�?            �F@       @7       8                 `�@1@      �?              @    �J@������������������������       �                     @      $@������������������������       �                      @      �?:       G                 �|Y=@�MI8d�?            �B@        ;       @                 ���@X�Cc�?             ,@      0@<       =                    5@���Q��?             @      @������������������������       �                     �?      �?>       ?                   �7@      �?             @      @������������������������       �                     @        ������������������������       �                     �?       @A       F                   �<@�<ݚ�?             "@     @B       C                   �8@      �?              @        ������������������������       �                     @        D       E                   @;@�q�q�?             @        ������������������������       �                     �?      @������������������������       �                      @      �?������������������������       �                     �?       @H       I                 ���@�nkK�?             7@        ������������������������       �                     @      �?J       M                 �|�=@      �?             0@       K       L                   @@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        O       V                 ���.@�q�q�?             (@       P       U                    �?      �?              @       Q       R                    �?r�q��?             @        ������������������������       �                     @        S       T                 �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X                       0�^I@Gq����?F           �@       Y       �                     @�"��c��?           P|@        Z       �                    �?z�7�Z�?\            @b@       [       t                 �|Y=@$��fF?�?L            @_@        \       a                    &@H�z�G�?             D@        ]       ^                    �?X�Cc�?             ,@        ������������������������       �                     @        _       `                   �7@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        b       k                   �;@�	j*D�?             :@       c       f                    �?�t����?             1@        d       e                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       h                    :@��S�ۿ?             .@       ������������������������       �        	             (@        i       j                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    �?�q�q�?             "@        ������������������������       �                     @        n       s                 `f�D@���Q��?             @       o       p                 `fF<@�q�q�?             @        ������������������������       �                     �?        q       r                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        u       �                   �*@ܻ�yX7�?1            @U@        v       }                   �>@��p\�?            �D@        w       x                    �?�r����?
             .@        ������������������������       �                     �?        y       |                 �|�=@@4և���?	             ,@       z       {                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ~                           �? ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �2@���|���?             F@ ,0,SOTO������������������������       �                     @ ,,1,0,3�       �                   @J@�z�G��?             D@le,30,0�       �                    �?�q�q�?             B@a Sophi�       �                    �?`�Q��?             9@ ussa, M������������������������       �                      @,"Jermy�       �                     �?��+7��?             7@, Mme. �       �                   �>@�z�G��?             4@,1,"Har�       �                 ��<:@�eP*L��?             &@ 
372,0,������������������������       �                      @ ,S
373,�       �                 X��B@�q�q�?             "@ ,S
374,������������������������       �                      @,C
375,0�       �                    H@և���X�?             @5,,S
37������������������������       �      �?             @ ,PC 176������������������������       �                     �? emale,2������������������������       �                     "@ male,27������������������������       �                     @e,20,0,�       �                    �?���|���?             &@ le,19,0�       �                   �E@�q�q�?             @,42,0,0������������������������       �                     @ ")",fem������������������������       �                      @ale,32,0������������������������       �                     @ exander������������������������       �                     @ 5,0,3,"�       �                    *@���N8�?             5@ 2,"Davi������������������������       �                      @ 87,0,3,�       �                    �?�S����?             3@,,S
388������������������������       �                     0@ ,"Sadli������������������������       �                     @mann, Mi�       �                    �?4����?�            0s@ Mr. Wil�       �                    �?      �?             L@ nsson, �       �                    @���B���?             :@afsson,�       �                    �?���}<S�?             7@Newell,�       �                 �|�9@      �?	             0@ 3,"Sand������������������������       �                     @4,0,2,P�       �                  ��@z�G�z�?             $@ 0,35005������������������������       �                      @50407,7������������������������       �                      @ 403,26,������������������������       �                     @400,1,2������������������������       �                     @ 12.65,,������������������������       �                     >@ 289,7.9�       �                    �?���w;�?�            `o@ S
403,0�       �                    �?�G�5��?)            @Q@
404,0,�       �                 ���1@b�2�tk�?             B@101279,�       �                 �|�<@��S���?             >@315096,�       �                 pf�@�q�q�?             2@ 21,,S
4������������������������       �                     @ 064,7.7�       �                   �2@z�G�z�?	             .@ 29106,1������������������������       �                     @21,0,0,�       �                    �?      �?             (@4133,25�       �                   �@�<ݚ�?             "@ 8958,,S�       �                 �&B@�q�q�?             @,1,1,"M�       �                   �7@      �?              @ ,2,"Cun������������������������       �                     �? 3,"Sund������������������������       �                     �? 5,,S
41������������������������       �                     �?0,0,3430������������������������       �                     @Christi�       �                 �!@�q�q�?             @ yyli Ka������������������������       �                     �?. Willi������������������������       �                      @. Cathar�       �                    �?�q�q�?	             (@ r. Stan�       �                   &@      �?             @id",mal������������������������       �                     @ ",male,������������������������       �                     �? t (Anna�       �                 ��Y.@      �?              @ 0,3,"Ro������������������������       �                     �?426,0,3������������������������       �                     @ 7,1,2,"������������������������       �                     @,0,2003,�       �                    :@�C��2(�?            �@@Louise �       �                   �6@@�0�!��?
             1@"Flynn,�       �                   �0@��S�ۿ?	             .@. Berk ������������������������       �                     "@,S
431,1�       �                    3@r�q��?             @ 0,11056������������������������       �                     �? nce Kat������������������������       �                     @ Charle������������������������       �                      @085,26,,������������������������       �                     0@O 2. 310�       �                 �?�@|)����?z            �f@ ,1,0,13�       �                    ?@@�)�n�?9            @U@,14,1,2�       �                    �?�\=lf�?-            �P@et ""Da�       �                 ���@ ������?)            �O@ ds, Mrs�       �                   �8@�����H�?             "@ 9,0,1,"�       �                   �4@z�G�z�?             @ 0,0,2,"������������������������       �                     �? 18723,1�       �                 �&b@      �?             @ d)",fem������������������������       �                     @ ",male,������������������������       �                     �?,male,25������������������������       �                     @female,������������������������       �        #             K@ Bernt",������������������������       �                     @ ton",ma�       �                 �&B@�����H�?             2@deleine������������������������       �                     (@r. Frede�       �                   �A@�q�q�?             @  Miss. �       �                   �@      �?             @ uchen, ������������������������       �                      @ ,0,2,"W������������������������       �                      @,0,3,"H������������������������       �                      @S
453,0�                          �?�*v��?A            @X@7.75,C1�       �                 @3�@ ��~���?<            �V@ ,89.104�       �                    �?X�Cc�?             ,@8.05,,S�       �                   �A@�	j*D�?             *@C
457,0�       �                   �:@"pc�
�?             &@ 8,S
458������������������������       �                     @64,51.86������������������������       ����Q��?             @C. 1353������������������������       �                      @ 0,7.75,������������������������       �                     �?E12,S
4�       �                    )@�KM�]�?4             S@ 63,0,1,������������������������       �                     �? ,"Milli�                          ?@���Lͩ�?3            �R@,"Maisn�                       �|�=@H�ՠ&��?$             K@ves, Mr�                          �?���C��?#            �J@S
467,0�                          �?�t����?!            �I@"Smart,�                       @3�!@(L���?            �E@,"Scanl�       �                 �|Y<@@�0�!��?             A@ Miss. �       �                 pf� @      �?             0@Keefe, �       �                 0S5 @"pc�
�?	             &@Luka",m�       �                   �3@�<ݚ�?             "@ ur (Ada�       �                   �1@      �?             @ Jerwan,������������������������       �                     �?H Basle������������������������       ��q�q�?             @ male,22������������������������       �                     @",male,,������������������������       �                      @ e,34,1,�       �                    8@���Q��?             @,1,0,34������������������������       �                     @ 0,0,350������������������������       �                      @,0,1,31�       �                 ��) @�����H�?
             2@,male,9������������������������       �                     .@ rchie""�                        pf� @�q�q�?             @ ",male,������������������������       �                      @ female,������������������������       �                     �?       ������������������������       �                     "@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @                                  @�q�q�?*            �L@       	      
                   �?���3�E�?%             J@       ������������������������       �                     @@                                 �?      �?             4@� t�q�                           �?�E��ӭ�?             2@                               �E@     ��?             0@                              x#J@�n_Y�K�?             *@        ������������������������       �                     @                                 �?      �?             $@        ������������������������       �                     �?                              `�iJ@X�<ݚ�?             "@        ������������������������       �                     @                              `f�N@�q�q�?             @                                7@      �?             @        ������������������������       �                     �?                                 A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @              !                   �?z�G�z�?             @                                  ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #      &                   �?h�����?             <@        $      %                  pE@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KM'KK��h]�Bp       0}@     �n@      .@     �@@      �?      =@              <@      �?      �?              �?      �?              ,@      @      $@              @      @       @               @      @              @       @             @|@     `j@     �z@     @j@     �M@     �P@      .@     �J@       @      A@       @      @       @                      @              <@      *@      3@      "@       @              �?      "@      @      @      @      @      @      @      @      @      @       @      @       @       @       @                       @              @       @              �?                      �?      �?              @              @      &@              @      @      @      @       @       @       @      �?       @      �?                       @      �?               @                       @      F@      *@     �B@       @      @       @      @                       @      ?@      @      "@      @       @      @      �?              �?      @              @      �?              @       @      @      �?      @               @      �?              �?       @                      �?      6@      �?      @              .@      �?      $@      �?      @      �?      @              @              @      @      @      �?      @      �?      @              �?      �?              �?      �?               @                      @     �v@      b@     �u@     �Z@     �W@      J@     @V@      B@      7@      1@      @      "@              @      @       @      �?       @      @              2@       @      .@       @      �?      �?              �?      �?              ,@      �?      (@               @      �?              �?       @              @      @              @      @       @      �?       @              �?      �?      �?              �?      �?               @             �P@      3@      C@      @      *@       @              �?      *@      �?      $@      �?      $@                      �?      @              9@      �?              �?      9@              <@      0@              @      <@      (@      8@      (@      1@       @               @      1@      @      ,@      @      @      @       @              @      @               @      @      @      @      @              �?      "@              @              @      @       @      @              @       @              @              @              @      0@       @              @      0@              0@      @             �o@      K@     �A@      5@      @      5@       @      5@       @      ,@              @       @       @       @                       @              @      @              >@             @k@     �@@      J@      1@      6@      ,@      0@      ,@      (@      @              @      (@      @      @              "@      @      @       @      �?       @      �?      �?              �?      �?                      �?      @               @      �?              �?       @              @       @      @      �?      @                      �?      �?      @      �?                      @      @              >@      @      ,@      @      ,@      �?      "@              @      �?              �?      @                       @      0@             �d@      0@     �T@      @     �P@      �?      O@      �?       @      �?      @      �?      �?              @      �?      @                      �?      @              K@              @              0@       @      (@              @       @       @       @               @       @               @              U@      *@     @S@      *@      "@      @      "@      @      "@       @      @              @       @               @              �?      Q@       @              �?      Q@      @     �G@      @     �G@      @     �F@      @     �B@      @      <@      @      (@      @      "@       @      @       @       @       @      �?              �?       @      @               @              @       @      @                       @      0@       @      .@              �?       @               @      �?              "@               @               @                      �?      5@              @              3@      C@      .@     �B@              @@      .@      @      *@      @      &@      @       @      @      @              @      @      �?              @      @              @      @       @       @       @      �?              �?       @               @      �?               @              @               @               @              @      �?      �?      �?              �?      �?              @              ;@      �?      �?      �?      �?                      �?      :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJؽ�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         P                     �?e�L��?�           8�@               3                    �?�G�z�?f             d@                                  �?���r
��?A            @X@  e n s                            �?�D����?             E@ \ g r                           @H@p�ݯ��?             C@     M@                        �|�;@�������?             >@      �?������������������������       �                     &@               	                    �?p�ݯ��?             3@     @������������������������       �                     $@�_4bQ  
                          �A@�<ݚ�?             "@^4bQ                          X�,@@����X�?             @[4bQ                          ��2>@r�q��?             @ ]4bQ  ������������������������       �                     �?�Y4bQ  ������������������������       �                     @0X4bQ  ������������������������       �                     �?�V4bQ  ������������������������       �                      @`U4bQ                          ��Z@      �?              @     �?������������������������       �                     @      �?������������������������       �                     �?      �?                        �\@      �?             @      �?������������������������       �                     �?      �?������������������������       �                     @      b@       *                 0�_J@N{�T6�?$            �K@     1@                           �?��.k���?             A@       @������������������������       �                     @      �?                        �|�<@���Q��?             >@        ������������������������       �                     @      @       )                    R@�q�q�?             ;@     �?       (                    L@�	j*D�?             :@              '                   �>@���Q��?             4@     �?                         �̌*@�q�q�?             (@      �?������������������������       �                      @        !       "                   �C@z�G�z�?             $@      (@������������������������       �                     @      @#       &                 `f�;@�q�q�?             @      @$       %                    H@z�G�z�?             @       ������������������������       �      �?             @      @������������������������       �                     �?      0@������������������������       �                     �?        ������������������������       �                      @      5@������������������������       �                     @        ������������������������       �                     �?        +       0                 03c@؇���X�?             5@     ,@,       -                    �?�IєX�?	             1@       ������������������������       �                     .@      �?.       /                    =@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?      @1       2                 ���f@      �?             @      @������������������������       �                      @      �?������������������������       �                      @        4       O                   �P@�<ݚ�?%            �O@     �?5       @                 ��Q@���*�?$             N@      �?6       7                    �?�q�q�?             2@        ������������������������       �                     @       @8       ?                    F@�eP*L��?             &@       9       :                    �?r�q��?             @      @������������������������       �                      @       @;       >                   @B@      �?             @     @<       =                   @K@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @        ������������������������       �                     �?       @������������������������       �                     @       @A       H                    �?���H��?             E@       B       G                    �?`Jj��?             ?@     C@C       D                    �?$�q-�?             :@     @������������������������       �        
             2@      @E       F                 ���^@      �?              @      @������������������������       �                     @       @������������������������       �                      @        ������������������������       �                     @      �?I       L                    �?���!pc�?             &@     �?J       K                 �U�X@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        M       N                 ��f`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Q       �                    �?�w�+`�?]           8�@       R       �                 Ь�#@�;�T<:�?           �z@       S       T                 ���@D�a�ў�?�            �p@        ������������������������       �                     <@        U       V                 ��@�.�PI�?�            �m@        ������������������������       �                     @        W       X                    /@P�z�?�            `m@        ������������������������       �                      @        Y       p                    �?F�|���?�             m@        Z       [                    �?Dc}h��?&             L@        ������������������������       �        	             *@        \       i                    �?�ʈD��?            �E@       ]       h                 �� @�LQ�1	�?             7@       ^       a                 ���@؇���X�?             5@        _       `                 �|�9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        b       g                 �|Y=@r�q��?	             (@        c       d                   @8@�q�q�?             @        ������������������������       �                     �?        e       f                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        j       k                 ���@P���Q�?             4@        ������������������������       �                     @        l       o                 X�I@      �?             0@       m       n                 ��(@��S�ۿ?             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        ������������������������       �                     �?        q       v                    �?$���?f             f@        r       u                   �@
;&����?             7@        s       t                   �A@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     &@        w       �                 �?�@�C��2(�?Z            @c@       x       y                 �|�<@����D��?5            @W@       ������������������������       �                     J@        z       �                   @@@������?            �D@       {       �                   �@�8��8��?             8@        |       �                 �&B@����X�?             @       }       ~                 ��@r�q��?             @        ������������������������       �                     @               �                 �|Y>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?  aQ  ������������������������       �        	             1@0aQ  ������������������������       �                     1@ �aQ  �       �                   �4@`��:�?%            �N@        �       �                   �0@�q�q�?
             .@        ������������������������       ����Q��?             @        �       �                 @3�@�z�G��?             $@        ������������������������       �                      @ aQ  �       �                 ��Y @      �?              @ �aQ  �       �                   �2@      �?             @        ������������������������       �                     �? �aQ  ������������������������       �                     @       ������������������������       �                     @       �       �                 @3�@*
;&���?             G@        �       �                   �A@      �?              @        ������������������������       �      �?             @ ,aQ  ������������������������       �      �?              @        �       �                    �?�˹�m��?             C@       �       �                 �|Y=@�8��8��?             B@        ������������������������       �                     "@ �aQ  �       �                 �|Y?@�����H�?             ;@vaQ  �       �                 ��) @r�q��?	             2@       ������������������������       �                     &@ aQ  �       �                 pf� @և���X�?             @        ������������������������       �                     @�aQ  ������������������������       �                     @        ������������������������       �                     "@ |aQ  ������������������������       �                      @        �       �                   �F@v�_���?e            �c@       �       �                   P,@�S��<�?Y            �a@ kaQ  �       �                    �?      �?$             N@        �       �                     @ 7���B�?             ;@       ������������������������       �                     4@ �aQ  �       �                    �?؇���X�?             @       �       �                 �[$@r�q��?             @        ������������������������       �                     @       �       �                 ��&@�q�q�?             @ �aQ  ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �%@<���D�?            �@@ ?aQ  ������������������������       �                     @        �       �                     @8�Z$���?             :@�aQ  �       �                 �|�<@�8��8��?             8@       ������������������������       �                     &@	aQ  �       �                 �|�=@8�Z$���?             *@ FaQ  ������������������������       �                      @       ������������������������       �                     &@        ������������������������       �                      @ �aQ  �       �                 pf�/@d�� z�?5            @T@ ?aQ  �       �                    1@      �?             0@ �aQ  �       �                   �-@      �?              @        ������������������������       �                     �?'aQ  ������������������������       �                     �?       ������������������������       �        
             ,@saQ  �       �                     @�4��?)            @P@       �       �                    �?؀�:M�?            �B@ �aQ  �       �                    �?      �?
             0@ �aQ  ������������������������       �                     @       �       �                    �?z�G�z�?             $@ 	aQ  ������������������������       �                     @aQ  �       �                   �;@����X�?             @ �aQ  ������������������������       �                     �? �aQ  �       �                   �E@r�q��?             @       ������������������������       �                     @       ������������������������       �                     �? �aQ  ������������������������       �                     5@ �aQ  �       �                 ���1@����X�?             <@        �       �                    �?      �?              @       ������������������������       �                     @ �aQ  ������������������������       �                     @ DaQ  �       �                    �?R���Q�?             4@ aQ  �       �                   �2@      �?              @        ������������������������       �                     @ �aQ  �       �                    �?���Q��?             @        ������������������������       �                      @3aQ  �       �                 �|�;@�q�q�?             @ �aQ  ������������������������       �                     �? 7aQ  ������������������������       �                      @       ������������������������       �                     (@        �       �                   �.@�IєX�?             1@       ������������������������       �        	             ,@       �       �                    5@�q�q�?             @ �aQ  ������������������������       �                     �? saQ  ������������������������       �                      @EaQ  �       �                     @X9����?U            �_@ �aQ  �       �                   �6@�������?             A@        ������������������������       �        
             .@ aQ  �       �                 ��J@�\��N��?             3@�aQ  �       �                    @���Q��?             .@�aQ  �       �                    �?X�Cc�?             ,@ �aQ  ������������������������       �                     @�aQ  ������������������������       �                     "@iaQ  ������������������������       �                     �?        ������������������������       �                     @ �aQ  �       �                    �?R�(��?=            @W@        �       �                 X��B@���y4F�?             3@eaQ  �       �                    @r�q��?             2@       �       �                    �?d}h���?             ,@       �       �                    3@r�q��?	             (@       �       �                    &@�q�q�?             @4aQ  ������������������������       �                     @       ������������������������       �                      @�aQ  ������������������������       �                     @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �? 6aQ  ������������������������       �                     @        ������������������������       �                     �?        �                       �̼6@^��4m�?0            �R@ aQ  �                       �̌5@�'�=z��?            �@@eaQ  �       �                   �*@*;L]n�?             >@        �       �                    (@�z�G��?             $@       ������������������������       �                     @�aQ  �       �                 xFT$@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @�aQ  �       �                    �?�z�G��?             4@       �       �                     @8�Z$���?	             *@aQ  �       �                    )@"pc�
�?             &@ �aQ  ������������������������       �                      @        ������������������������       �                     "@       ������������������������       �                      @paQ  �       �                 @33/@և���X�?             @        ������������������������       �                     �? �aQ  �                           �?�q�q�?             @        ������������������������       �                     @                                 +@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        ������������������������       �                     @              
                   �?��p\�?            �D@              	                  @C@�t����?
             1@                                �B@      �?              @       ������������������������       �                     @        ������������������������       �                      @       ������������������������       �                     "@                              ��p@@ �q�q�?             8@ � ��q�                       ��T?@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        
             *@        �t�b��     h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@      J@      [@      C@     �M@      1@      9@      ,@      8@      @      7@              &@      @      (@              $@      @       @      @       @      @      �?              �?      @                      �?       @              @      �?      @                      �?      @      �?              �?      @              5@      A@      2@      0@              @      2@      (@              @      2@      "@      2@       @      (@       @      @       @       @               @       @              @       @      @      �?      @      �?      @              �?      �?               @              @                      �?      @      2@      �?      0@              .@      �?      �?              �?      �?               @       @       @                       @      ,@     �H@      &@     �H@      @      (@              @      @      @      �?      @               @      �?      @      �?       @      �?                       @              �?      @              @     �B@       @      =@       @      8@              2@       @      @              @       @                      @      @       @      �?      @              @      �?               @       @       @                       @      @             px@      d@     0t@     @Y@     `k@     �G@      <@             �g@     �G@              @     �g@      F@               @     �g@      E@     �C@      1@              *@     �C@      @      4@      @      2@      @       @      �?              �?       @              $@       @      �?       @              �?      �?      �?      �?                      �?      "@               @              3@      �?      @              .@      �?      ,@      �?      (@      �?       @              �?              c@      9@      (@      &@      �?      &@              &@      �?              &@             �a@      ,@     �V@       @      J@             �C@       @      6@       @      @       @      @      �?      @               @      �?      �?      �?      �?                      �?      1@              1@             �H@      (@      $@      @      @       @      @      @               @      @      �?      @      �?              �?      @              @             �C@      @      @      @      @      @      �?      �?     �A@      @     �@@      @      "@              8@      @      .@      @      &@              @      @              @      @              "@               @              Z@      K@      V@     �J@      >@      >@      �?      :@              4@      �?      @      �?      @              @      �?       @      �?                       @              �?      =@      @      @              6@      @      6@       @      &@              &@       @               @      &@                       @      M@      7@      .@      �?      �?      �?      �?                      �?      ,@             �E@      6@      7@      ,@       @      ,@              @       @       @              @       @      @      �?              �?      @              @      �?              5@              4@       @      @      @              @      @              1@      @      @      @      @               @      @               @       @      �?              �?       @              (@              0@      �?      ,@               @      �?              �?       @              Q@     �M@      "@      9@              .@      "@      $@      "@      @      "@      @              @      "@                      �?              @     �M@      A@      @      .@      @      .@      @      &@       @      $@       @      @              @       @                      @      �?      �?              �?      �?                      @      �?             �K@      3@      1@      0@      1@      *@      @      @              @      @       @      @                       @      ,@      @      &@       @      "@       @               @      "@               @              @      @      �?               @      @              @       @      �?              �?       @                      @      C@      @      .@       @      @       @      @                       @      "@              7@      �?      $@      �?      $@                      �?      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX��vhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@A         d                    �?e�L��?�           8�@               _                    @<�T]���?�            �o@     @       \                    @Q��"�?�            `m@      @       G                 �|�=@��^���?�             m@    �M@                           !@ܱ#_��?\            `b@        ������������������������       �                     ,@      @                           '@���c�?T            �`@      �?������������������������       �                     @       @	                            @:�����?R            �_@        
                           �?���J��?"            �I@      @������������������������       �                     4@      �?                           �?�g�y��?             ?@                                  9@P���Q�?             4@      =@                           �?      �?             @                                 �'@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      2@������������������������       �                      @      @������������������������       �                     0@        ������������������������       �                     &@               :                    �?���=A�?0             S@              %                 @� @     ��?)             P@      @                          �6@��s����?             E@      @������������������������       �        
             4@      �?                          �9@���|���?             6@      �?                        pf�@      �?             @        ������������������������       �                     �?      �?������������������������       �                     @                                   ;@�E��ӭ�?             2@      &@������������������������       �                      @       @       $                    �?     ��?             0@      @        #                 ���@d}h���?	             ,@      �?!       "                 �Y�@���Q��?             @        ������������������������       �                      @      @������������������������       �                     @      �?������������������������       �                     "@      @������������������������       �                      @      @&       1                    �?8�A�0��?             6@        '       (                   �,@      �?             (@        ������������������������       �                      @      >@)       0                    �?�z�G��?             $@     @*       /                  S�-@�q�q�?             "@      @+       .                 �|Y6@���Q��?             @     @,       -                   �-@�q�q�?             @       @������������������������       �                     �?      �?������������������������       �                      @        ������������������������       �                      @      @������������������������       �                     @        ������������������������       �                     �?        2       9                 �|�:@���Q��?	             $@       3       8                    �?؇���X�?             @     @4       5                  �#@      �?             @        ������������������������       �                      @      �?6       7                 �[$@      �?              @      9@������������������������       �                     �?      @������������������������       �                     �?      @������������������������       �                     @      &@������������������������       �                     @        ;       @                   �6@�q�q�?             (@        <       ?                   �3@z�G�z�?             @     0@=       >                    �?      �?             @       @������������������������       �                     @       @������������������������       �                     �?        ������������������������       �                     �?      @A       B                 �|�:@և���X�?             @      �?������������������������       �                      @ 6aQ  C       D                    �?z�G�z�?             @ �aQ  ������������������������       �                      @ �aQ  E       F                    �?�q�q�?             @      �?������������������������       �                     �?PaQ  ������������������������       �                      @       @H       W                    �?�̨�`<�?8            @U@"aQ  I       J                   @B@؇���X�?%             L@"aQ  ������������������������       �                     ;@ (aQ  K       V                 83'E@�c�Α�?             =@�aQ  L       O                     �?      �?	             0@ �aQ  M       N                    �?؇���X�?             @ -aQ  ������������������������       �                     �? �aQ  ������������������������       �                     @ aQ  P       U                   �+@�<ݚ�?             "@       Q       T                     @�q�q�?             @aQ  R       S                    D@���Q��?             @ �aQ  ������������������������       �                     @ aQ  ������������������������       �                      @�aQ  ������������������������       �                     �? haQ  ������������������������       �                     @�LaQ  ������������������������       �                     *@ �aQ  X       Y                     @XB���?             =@^aQ  ������������������������       �                     7@ aQ  Z       [                    C@r�q��?             @ �aQ  ������������������������       �                     @aQ  ������������������������       �                     �? aQ  ]       ^                 ��T?@�q�q�?             @�aQ  ������������������������       �                      @ aQ  ������������������������       �                     �? BaQ  `       a                      @�t����?             1@ �aQ  ������������������������       �                     @        b       c                 �|Y?@$�q-�?
             *@aQ  ������������������������       �        	             (@        ������������������������       �                     �?       e       �                 ��K.@�#2����?"           �|@�aQ  f       w                    �?�]l*7��?�            0r@ �aQ  g       h                   �6@>���Rp�?             M@ �aQ  ������������������������       �                     "@ �aQ  i       n                 �|Y=@ i���t�?            �H@ KaQ  j       m                    �?      �?             (@       k       l                   �<@�q�q�?             "@�aQ  ������������������������       �                     @ =aQ  ������������������������       �                     @aaQ  ������������������������       �                     @ aQ  o       p                 ���@@-�_ .�?            �B@ %aQ  ������������������������       �                     .@ &aQ  q       r                     @�C��2(�?             6@ �aQ  ������������������������       �                     @ �aQ  s       v                 �|�=@�����H�?	             2@       t       u                   @@"pc�
�?             &@       ������������������������       �����X�?             @       ������������������������       �                     @ �aQ  ������������������������       �                     @�aQ  x       �                    �?`�q��־?�             m@�aQ  y       �                 ���"@ �Cc��?�             l@�aQ  z       �                 ��@�1��?o            �e@        {       |                     @��v$���?*            �N@ �aQ  ������������������������       �                     $@aQ  }       �                 ���@���J��?#            �I@ )aQ  ~                        ���@�IєX�?
             1@�aQ  ������������������������       �        	             0@9aQ  ������������������������       �                     �? �aQ  ������������������������       �                     A@ ,4,4,2,�       �                    �?�h����?E             \@0,34706�       �                   �3@ ѯ��?B            �Z@ ,2678,1�       �                   �1@��2(&�?             6@ ,1,PC 1������������������������       �                     &@Lilian H�       �                 �?�@���!pc�?             &@  (Leah ������������������������       �                     @ George �       �                 ��Y @���Q��?             @
858,1,�       �                   �2@      �?             @ 
859,1,������������������������       �                      @666,19.������������������������       �      �?              @ ,C
861,������������������������       �                     �?,,S
862,�       �                 �|Y=@@�)�n�?6            @U@ ,S
863,������������������������       �                    �B@,female�       �                   @@@      �?             H@Edith "�       �                    ?@�#-���?            �A@. John �       �                 �|�=@@4և���?             <@(Karoli�       �                  sW@HP�s��?             9@ ss. Asu������������������������       �      �?             @ ebling,������������������������       �                     5@ ,A24,S
������������������������       �                     @.5,,S
87�       �                 P�@؇���X�?             @ ,11.133������������������������       �                     �?58,,S
87������������������������       �                     @ female,������������������������       �                     *@ lof",ma������������������������       �                     @Mr. Vict�       �                   @B@�t����?$            �I@ (Hanna�       �                   �@@R���Q�?             D@ Miss. �       �                     @�ݜ�?            �C@3,"Gust�       �                    5@���7�?             6@ ,0,3,"P�       �                   �2@z�G�z�?             @ ,"Lalef������������������������       �                      @ , Mrs. ������������������������       ��q�q�?             @ 1583,C5������������������������       �                     1@",femal�       �                 `�X#@������?             1@3,0,0,3�       �                   �<@�	j*D�?             *@ male,22������������������������       �                     @ es",mal�       �                 �|Y=@X�<ݚ�?             "@ Henry J������������������������       �                      @ . Willi�       �                 �|�=@����X�?             @ 0,2,"Mo������������������������       �                     @ aham, M�       �                   �?@      �?             @ 3,"John������������������������       �                      @  6607,2������������������������       �                      @ 9,30,C1������������������������       �                     @75,,Q
  ������������������������       �                     �?       ������������������������       �                     &@       �       �                    �?�<ݚ�?             "@        ������������������������       �                      @       �       �                    �?����X�?             @       �       �                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@      �?l             e@       �       �                   @A@�Sb(�	�?D             [@       �       �                 `�/@�Y|���?A            �Y@        ������������������������       �                     @       �       �                    @�D��??            �X@       �       �                    �?^H���+�?3            �R@       �       �                    �?�Gi����?            �B@       �       �                    �?���|���?            �@@        �       �                      @�q�q�?             "@       �       �                 �|Y<@����X�?             @        �       �                    9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �?@      �?             8@       �       �                 `f�D@����X�?             5@       �       �                     �?��
ц��?	             *@       �       �                   �<@�q�q�?             "@        ������������������������       �                      @       �       �                 `fF<@և���X�?             @        ������������������������       �                      @        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 h"_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?V������?            �B@        �       �                    �?�<ݚ�?             "@       �       �                    ;@      �?              @       �       �                    �?���Q��?             @       �       �                 8�T@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?       �       �                    )@��X��?             <@        ������������������������       �                     @        �       �                 `fFJ@�����?             5@       ������������������������       �        
             .@        �       �                     �?�q�q�?             @       �       �                    7@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     8@        �       �                     �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?�?�P�a�?(             N@       �       �                    H@r�q��?             E@       �       �                    �?`2U0*��?             9@       �       �                    �?      �?	             0@        ������������������������       �                     �?        �       �                   �F@��S�ۿ?             .@        �       �                 `fF:@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     "@       �                       �5L@ҳ�wY;�?             1@       �                        i?@������?
             .@       �       �                 `fF:@���|���?             &@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?                                 L@և���X�?             @        ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �t�bh�h*h-K ��h/��R�(KMKK��h]�BP       �{@     �p@     �K@     �h@     �E@      h@     �D@     �g@      @@     �\@              ,@      @@     @Y@      @              :@     @Y@      �?      I@              4@      �?      >@      �?      3@      �?      @      �?      �?              �?      �?                       @              0@              &@      9@     �I@      1@     �G@       @      A@              4@       @      ,@      @      �?              �?      @              @      *@               @      @      &@      @      &@      @       @               @      @                      "@       @              "@      *@      @      "@               @      @      @      @      @      @       @      �?       @      �?                       @       @                      @              �?      @      @      @      �?      @      �?       @              �?      �?              �?      �?              @                      @       @      @      @      �?      @      �?      @                      �?      �?              @      @               @      @      �?       @               @      �?              �?       @              "@      S@       @      H@              ;@       @      5@       @       @      �?      @      �?                      @      @       @      @       @      @       @      @                       @      �?              @                      *@      �?      <@              7@      �?      @              @      �?               @      �?       @                      �?      (@      @              @      (@      �?      (@                      �?     @x@     �Q@     `p@      =@      F@      ,@              "@      F@      @      "@      @      @      @      @                      @      @             �A@       @      .@              4@       @      @              0@       @      "@       @      @       @      @              @             @k@      .@     `j@      *@     �d@      @      N@      �?      $@              I@      �?      0@      �?      0@                      �?      A@             �Z@      @     @Y@      @      3@      @      &@               @      @      @               @      @      �?      @               @      �?      �?      �?             �T@      @     �B@             �F@      @      @@      @      :@       @      7@       @       @       @      5@              @              @      �?              �?      @              *@              @             �F@      @      A@      @      A@      @      5@      �?      @      �?       @               @      �?      1@              *@      @      "@      @      @              @      @               @      @       @      @               @       @               @       @              @                      �?      &@              @       @       @              @       @      @       @               @      @               @             �_@      E@     @R@     �A@      R@      ?@              @      R@      :@      H@      :@      6@      .@      5@      (@      @      @      @       @      �?       @      �?                       @      @              �?      �?      �?                      �?      .@      "@      .@      @      @      @      @      @               @      @      @       @              �?      @      �?                      @      @               @                      @      �?      @              @      �?              :@      &@      @       @      @       @      @       @       @       @               @       @              �?              @              �?              3@      "@              @      3@       @      .@              @       @      �?       @      �?                       @      @              8@              �?      @              @      �?             �J@      @     �A@      @      8@      �?      .@      �?      �?              ,@      �?      @      �?      @               @      �?      "@              "@              &@      @      &@      @      @      @      @              @      @      �?              @      @              @      @              @                       @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���EhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         r                     @�����?�           8�@                                   �?yÏP�?�            �t@      �?                        03�<@@+K&:~�?[             c@      @                           �?Xny��?(            �N@                                 �H@>A�F<�?             C@     M@                           �?�t����?             A@     �?                          @B@�nkK�?             7@       ������������������������       �                     2@     @	       
                   �,@z�G�z�?             @        ������������������������       �                     �?      @������������������������       �                     @      �?                           �?���!pc�?             &@        ������������������������       �                     �?      =@                          �;@�z�G��?             $@                                  �7@�q�q�?             @        ������������������������       �                      @      @������������������������       �                     �?      2@                           D@؇���X�?             @     @������������������������       �                     @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                      @      @                          �J@      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      �?������������������������       �                     7@        ������������������������       �        3            �V@      �?       =                    �?:���١�?p             f@               8                     �?�[�IJ�?            �G@     &@       5                    �?      �?             C@      @                         ��";@��>4և�?             <@       @������������������������       �                      @      �?!       4                 �̾w@$��m��?             :@     @"       '                 �|Y<@`�Q��?             9@       @#       &                    �?      �?              @      @$       %                  �}S@և���X�?             @     $@������������������������       �                     @      @������������������������       �                     @       @������������������������       �                     �?      @(       3                    �?@�0�!��?             1@     :@)       2                 p�i@@�θ�?	             *@      @*       /                   �A@և���X�?             @     �?+       ,                 ���<@      �?             @      &@������������������������       �                      @      @-       .                 ��2>@      �?              @       @������������������������       �                     �?     �?������������������������       �                     �?      @0       1                  �>@�q�q�?             @       @������������������������       �                     �?       @������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     @      P@������������������������       �                     �?     @6       7                 ��>Y@z�G�z�?             $@      @������������������������       �                      @    �J@������������������������       �                      @      $@9       :                    �?�����H�?             "@     �?������������������������       �                     @        ;       <                 pV�C@      �?              @      0@������������������������       �                     �?      @������������������������       �                     �?      �?>       m                    �?
�e4���?Q             `@     @?       Z                     �?d�X^_�?I            �\@        @       O                    B@H.�!���?!             I@       @A       N                 `f�D@�LQ�1	�?             7@      @B       C                 ��I*@��S���?
             .@        ������������������������       �                     @        D       E                   �<@z�G�z�?             $@        ������������������������       �                     @        F       M                   @>@����X�?             @       G       L                 �|�?@���Q��?             @       H       I                 �|Y=@�q�q�?             @        ������������������������       �                     �?        J       K                 `fF<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        P       Y                 ���[@�����H�?             ;@       Q       X                    �?$�q-�?             :@       R       W                 `f�;@�C��2(�?             6@       S       V                   �K@r�q��?             (@        T       U                 ��:@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     �?        [       l                    �?P�2E��?(            @P@       \       k                   �*@�X�<ݺ?              K@       ]       ^                   �(@$�q-�?            �C@        ������������������������       �        	             ,@        _       `                 �|�<@H%u��?             9@        ������������������������       �                     "@        a       b                 �|�=@     ��?             0@        ������������������������       �                     �?        c       j                   �F@�r����?
             .@       d       i                   @D@z�G�z�?             $@       e       f                    @@�����H�?             "@        ������������������������       �                     @        g       h                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     &@        n       o                    :@X�Cc�?             ,@        ������������������������       �                     @        p       q                    5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        s                          @l���`��?�            �w@       t       �                    �?B�>�;Q�?�            �w@       u       �                    �?C؇eY�?�            �p@        v                        P��@�ucQ?-�?3            @U@        w       ~                 ���@      �?             8@       x       y                 03S@z�G�z�?
             .@        ������������������������       �                     �?        z       {                   �7@d}h���?	             ,@        ������������������������       �                      @        |       }                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     "@        �       �                    �?��7��?#            �N@       �       �                 �|Y=@\X��t�?             G@ 910,15.�       �                    �?     ��?	             0@ 58,,S
6�       �                   �2@      �?             @ 0.5,,S
������������������������       �                     �?rgue)",������������������������       �                     @ iss. El�       �                    �?r�q��?             (@,"Ander������������������������       �                      @ale,39,�       �                    ;@      �?             @ ,,0,0,S������������������������       �                      @  Jane",������������������������       �                      @ e,,0,0,�       �                    �?�������?             >@ male,35������������������������       �                     @ 24,1,2,�       �                 @a'@8����?             7@1,1,347�       �                 `�j@�q�q�?             5@K Stanl�       �                 X��A@�z�G��?             4@ss. Mar�       �                 �;@�����?             3@r. Lawr�       �                 03@�q�q�?             2@oni",ma�       �                 ��@�t����?             1@ son Jr"�       �                    �?      �?              @ d",male������������������������       �                     �? ard",ma������������������������       �                     �?  ""Dai"�       �                 ���@������?	             .@ ck",mal������������������������       �                     �? les Leo�       �                    �?����X�?             ,@  Gretch������������������������       �                     @ndyeff,������������������������       �                     $@nnell, ������������������������       �                     �?rth, Mr������������������������       �                     �? ,3,"Lun������������������������       �                     �? 3,1,1,"������������������������       �                     �? 34,0,1,������������������������       �                      @ ,0,3,"S�       �                    �?z�G�z�?             .@ avis, M�       �                    &@      �?              @ Mr. Ant������������������������       �                      @,"Colly������������������������       �                     @ Panula,�       �                 ���&@؇���X�?             @ .6875,,������������������������       �                     @6.1,,S
�       �                 �|Y=@      �?             @ 2,,S
64������������������������       �                     �? B35,C
6������������������������       �                     @ 8,27.9,�       �                   �0@X��Oԣ�?t            @g@ 5,1,3,"������������������������       �                     @ 46,1,1,�       �                    �?�8��8��?o            �f@ D33,C
6�       �                 ���@�q�q�?
             .@ 48,1,1,������������������������       �                     �?5.5,A26�       �                 �|�;@����X�?	             ,@.55,,S
�       �                   �9@���|���?             &@A. 2314�       �                    8@�<ݚ�?             "@958,,S
�       �                   �6@����X�?             @653,0,3�       �                  �#@r�q��?             @,,S
654������������������������       �                     @ ,7.8292������������������������       �                     �?0,36522������������������������       �                     �? ,S.O.C.������������������������       �                      @349223,������������������������       �                      @32,1,1,������������������������       �                     @ e,23,0,�       �                 �?�@�FVQ&�?e            �d@ 8,0,2,3�       �                 �|Y=@`<)�+�?1            @S@",male,�       �                   �8@p���?             I@e,40,0,�       �                   �7@ ��WV�?             :@,47,0,0������������������������       �                     7@0,34921�       �                 `fF@�q�q�?             @ ,1,0,ST������������������������       �                     �? e,32,2,������������������������       �                      @on",mal������������������������       �                     8@",male,�       �                 �|Y>@�>����?             ;@ 0,A/5 3�       �                  sW@�t����?
             1@ mmins W�       �                 ��,@�q�q�?             @ Thomas ������������������������       �                     @ ,29750,������������������������       ��q�q�?             @2750,52������������������������       �                     &@C.A. 24������������������������       �        
             $@ 44270,1�       �                   �3@`���i��?4             V@ 6,0,,S
�       �                   �1@�θ�?             *@ 12,7.77������������������������       �                      @ 0,34282�       �                 `�8"@���!pc�?             &@,4138,9�       �                   �2@և���X�?             @ ",femal������������������������       �                     �? ke Mart������������������������       ��q�q�?             @,"Peter������������������������       �                     @ sab, Mr�       �                   �:@Х-��ٹ?-            �R@ vigen, ������������������������       �                     <@dwin, M�       �                   �;@dP-���?             �G@ rown, M������������������������       �                     �? 2,"Laro�       �                 @3�@���.�6�?             G@ 2123,41�       �                   �?@�q�q�?             @ 101295,������������������������       �                     �?,10.170������������������������       �                      @ 0,35003�       �                 ��) @ �#�Ѵ�?            �E@ emale,1������������������������       �                     7@ n",male�       �                 �|�>@ףp=
�?             4@e,4,0,1�       �                 pf� @r�q��?
             (@ 56.4958������������������������       �                     �?695,0,1�       �                    (@�C��2(�?	             &@ hapman,�       �                 �|Y=@z�G�z�?             @ elly, M�       �                 ���"@      �?              @ ss. Kat������������������������       �                     �?ayer, M������������������������       �                     �?,"Humbl������������������������       �                     @ .65,F G������������������������       �                     @Force)"������������������������       �                      @thorne,�                          �?������?L             [@03,0,3,�       �                    �?�BE����?)             O@ ,0,3,"G�       �                    �?      �?             $@,"Hanse�       �                    �?X�<ݚ�?             "@"Morley�       �                  S�-@����X�?             @ 50655,2�       �                 03�)@�q�q�?             @ 0,0,223������������������������       �                     �? ale,42,������������������������       �                      @ ,female������������������������       �                     @  Gonios������������������������       �                      @,"Mayne,������������������������       �                     �? ,0,PC 1�       �                    �?�	j*D�?!             J@,113028�       �                   �3@�P�*�?             ?@ 1,0,199������������������������       �                     @ ,0,0,75�       �                 �|Y=@�q�q�?             ;@ 250647,������������������������       �                     *@ ",male,�       �                 03�1@X�Cc�?             ,@ e Louis�       �                 ���.@ףp=
�?             $@ Miss. E������������������������       �                     �? 19,0,3,������������������������       �                     "@hnson, ������������������������       �                     @,"Harper�                          �?؇���X�?             5@722,0,3�                          �?�KM�]�?             3@
723,0,�                        ��y'@�8��8��?	             (@ 724,0,2�       �                 P�@z�G�z�?             @,1,"Cha������������������������       �                     @ 726,0,3������������������������       �                     �? ,2,"Ren������������������������       �                     @                                $@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?*
;&���?#             G@        	                      ��*4@��<b���?             7@        
                        �1@      �?             @        ������������������������       �                      @�� 1�q�                          @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @�KM�]�?             3@                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@                                 �?���}<S�?             7@       ������������������������       �                     *@                                 @z�G�z�?             $@                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �a@     �g@      @      b@      @      K@      @      ?@      @      >@      �?      6@              2@      �?      @      �?                      @      @       @              �?      @      @       @      �?       @                      �?      �?      @              @      �?              @      �?       @              �?      �?              �?      �?                      7@             �V@     �`@     �E@      ;@      4@      3@      3@      1@      &@               @      1@      "@      1@       @      @      @      @      @              @      @                      �?      ,@      @      $@      @      @      @      @      �?       @              �?      �?              �?      �?              �?       @      �?                       @      @              @                      �?       @       @               @       @               @      �?      @              �?      �?              �?      �?             �Z@      7@     @Y@      ,@     �C@      &@      .@       @      @       @      @               @       @              @       @      @       @      @       @      �?      �?              �?      �?      �?                      �?               @               @       @              8@      @      8@       @      4@       @      $@       @      @       @      @                       @      @              $@              @                      �?      O@      @     �I@      @      B@      @      ,@              6@      @      "@              *@      @              �?      *@       @       @       @       @      �?      @              @      �?       @      �?      @                      �?      @              .@              &@              @      "@              @      @       @               @      @              s@     @S@      s@     �R@      l@     �G@     �M@      :@      5@      @      (@      @      �?              &@      @               @      &@      �?              �?      &@              "@              C@      7@      :@      4@      @      *@      �?      @      �?                      @       @      $@               @       @       @       @                       @      7@      @      @              0@      @      ,@      @      ,@      @      *@      @      (@      @      (@      @      �?      �?              �?      �?              &@      @      �?              $@      @              @      $@                      �?      �?              �?                      �?       @              (@      @      @       @               @      @              @      �?      @              @      �?              �?      @             �d@      5@              @     �d@      .@      $@      @              �?      $@      @      @      @      @       @      @       @      @      �?      @                      �?              �?       @                       @      @             `c@      $@     �R@      @     �H@      �?      9@      �?      7@               @      �?              �?       @              8@              9@       @      .@       @      @       @      @              �?       @      &@              $@             @T@      @      $@      @       @               @      @      @      @              �?      @       @      @             �Q@      @      <@             �E@      @              �?     �E@      @       @      �?              �?       @             �D@       @      7@              2@       @      $@       @              �?      $@      �?      @      �?      �?      �?      �?                      �?      @              @               @              T@      <@     �D@      5@      @      @      @      @       @      @       @      �?              �?       @                      @       @              �?              B@      0@      2@      *@              @      2@      "@      *@              @      "@      �?      "@      �?                      "@      @              2@      @      1@       @      &@      �?      @      �?      @                      �?      @              @      �?              �?      @              �?      �?              �?      �?             �C@      @      2@      @      �?      @               @      �?      �?      �?                      �?      1@       @      �?       @      �?                       @      0@              5@       @      *@               @       @      �?       @               @      �?              @               @       @      �?              �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:9)bhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         �                     @e�L��?�           8�@      K@       Y                     �?x@����?�            �u@               P                   �J@���(�_�?k            �e@     @                        `V�9@�ӭ�a�?Y             b@      �?������������������������       �                     @                                  �7@�:���?T             a@      @������������������������       �                     3@      �?       %                   �?@�k��(A�?I            �]@       @	                         x;K@Fx$(�?             I@��XQ  
                          �<@|��?���?             ;@ ��XQ  ������������������������       �                      @���XQ                            �>@�����?             3@pDYQ                          �|Y=@���Q��?	             .@ ��XQ  ������������������������       �                      @\�XQ                            �<@��
ц��?             *@ ��XQ  ������������������������       �                     @ ��XQ                            @D@���Q��?             $@      @������������������������       �                     @      .@                          �I@z�G�z�?             @      (@������������������������       �                      @      �?                           �?�q�q�?             @      @������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               "                    �?��+7��?             7@     @                           �?�t����?             1@       ������������������������       �                     (@      �?                        `f�N@���Q��?             @      @������������������������       �                      @     �D@       !                    �?�q�q�?             @     @                          �}S@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                     �?       @#       $                    �?�q�q�?             @       ������������������������       �                     @      @������������������������       �                      @      �?&       E                 x5Q@�M���?*             Q@     @'       D                 0��M@ҳ�wY;�?             A@       (       1                 ���;@¦	^_�?             ?@      @)       *                 03k:@8�Z$���?             *@      �?������������������������       �                     @        +       ,                    �?z�G�z�?             $@      @������������������������       �                     �?       @-       .                   �C@�<ݚ�?             "@      �?������������������������       �                     @        /       0                    H@�q�q�?             @     �?������������������������       �      �?             @        ������������������������       �                      @       @2       5                    �?b�2�tk�?             2@        3       4                 ��A@      �?              @      @������������������������       �                      @        ������������������������       �                     @      �?6       ;                    �?      �?             $@        7       :                    �?      �?             @      @8       9                    C@�q�q�?             @      �?������������������������       �                      @        ������������������������       �                     �?      @������������������������       �                     �?      �?<       =                   �C@      �?             @        ������������������������       �                     �?      "@>       A                    �?���Q��?             @        ?       @                   @A@      �?              @       @������������������������       �                     �?      �?������������������������       �                     �?      &@B       C                 �K@�q�q�?             @      �?������������������������       �                      @        ������������������������       �                     �?      6@������������������������       �                     @      @F       G                    �?l��\��?             A@       ������������������������       �        
             0@        H       I                    �?r�q��?	             2@        ������������������������       �                      @        J       O                    �?�z�G��?             $@       K       N                 Ј�U@      �?              @        L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                 �U'Q@ܷ��?��?             =@       ������������������������       �                     6@        S       T                    �?և���X�?             @        ������������������������       �                      @        U       V                   �K@z�G�z�?             @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �1@և���X�?k            �e@        [       \                    �?�}�+r��?             3@       ������������������������       �                     ,@        ]       ^                    #@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �                    L@����3��?_            �c@       a       |                    �?Fx$(�?Y            �b@        b       {                    :@��ϭ�*�?'             M@       c       d                    �?�����H�?            �F@        ������������������������       �                     @        e       z                    �?,���i�?            �D@       f       s                    �?6YE�t�?            �@@       g       j                   �9@�C��2(�?             6@        h       i                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �'@�}�+r��?             3@        ������������������������       �                     @        m       r                   �,@�8��8��?             (@       n       o                    B@�����H�?             "@       ������������������������       �                     @        p       q                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       y                   �E@���!pc�?             &@       u       x                   �;@�����H�?             "@        v       w                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        }       ~                 �|Y=@�nkK�?2             W@        ������������������������       �                     A@               �                   �*@ 	��p�?!             M@       �       �                    �?(N:!���?            �A@        ������������������������       �                     @, Mr. N�       �                 �|�=@      �?             @@ �GbQ  �       �                    @�q�q�?             "@�GbQ  ������������������������       �                     @ GbQ  ������������������������       �                     @ McMahon�       �                   @D@�nkK�?             7@r. Frid������������������������       �                     &@ Miss. A�       �                 `f�)@�8��8��?             (@ r. Joha������������������������       �                      @9GbQ  �       �                   �F@ףp=
�?             $@ GbQ  ������������������������       ��q�q�?             @ns, Mrs.������������������������       �                     @GbQ  ������������������������       �                     7@ )",fema������������������������       �                     @ayden",�       �                    @��,?S�?�            �v@ ,male,2�       �                    @$��m��?             :@ en Mony������������������������       �                     &@��GbQ  �       �                    @���Q��?             .@n, Mr. ������������������������       �                     @. Victo�       �                    �?      �?              @ Joseph ������������������������       �                      @ �FbQ  �       �                 ��T?@�q�q�?             @ �GbQ  ������������������������       �                      @O2. 310������������������������       �                     @�$GbQ  �       �                    �?�B���?�            u@ 31945,1�       �                   @C@     ��?=             X@GbQ  �       �                    �?V�K/��?5            �S@ nnerstr�       �                    �?���B���?             :@aGbQ  �       �                    �?P���Q�?             4@ 2,"Navr�       �                 ���,@      �?             @080,26,������������������������       �                     @��GbQ  ������������������������       �                     �? 0,S.O.P������������������������       �                     0@e)",fem�       �                 `�@1@�q�q�?             @�FbQ  �       �                    �?z�G�z�?             @  Blyler������������������������       �                      @ Martin"�       �                 �|Y=@�q�q�?             @ rles Du������������������������       �                     �? <8bQ  ������������������������       �                      @"Corn, M������������������������       �                     �? iljanic�       �                   @A@Fmq��?             �J@ter. Th�       �                   @1@���Q �?            �H@�GbQ  �       �                    �?)O���?             B@ James �       �                   �5@8�A�0��?             6@ �FbQ  �       �                   �3@؇���X�?             @47068,7�       �                   !@      �?              @ .GbQ  ������������������������       �                     �?�GbQ  ������������������������       �                     �?kie""",������������������������       �                     @h Marth�       �                 �|�=@��S���?             .@�FbQ  �       �                 ��&@�n_Y�K�?
             *@�GbQ  �       �                    ;@���!pc�?             &@�0bQ  �       �                 03�!@և���X�?             @an der �       �                   �7@      �?             @ �GbQ  ������������������������       �                      @son, Mi�       �                 pff@      �?              @ �GbQ  ������������������������       �                     �? ,,S
175������������������������       �                     �?58bQ  ������������������������       �                     @ ?8bQ  ������������������������       �                     @7,,S
17������������������������       �                      @-GbQ  ������������������������       �                      @ =GbQ  �       �                    �?����X�?             ,@�FbQ  �       �                    �?�θ�?             *@�FbQ  �       �                 ���)@�q�q�?             "@ 3,"Aspl������������������������       �                     @ 875,,S
�       �                 �|�;@      �?             @ �6bQ  ������������������������       �                     �?��FbQ  ������������������������       �                     @ 7,50,A3������������������������       �                     @frey)",������������������������       �                     �? 5bQ  ������������������������       �        	             *@0�GbQ  ������������������������       �                     @ <GbQ  ������������������������       �                     1@ Rosa)",�                          �?P�_��I�?�             n@
GbQ  �       �                    �?      �?�             l@ Christi�       �                 �=/@�<ݚ�?$             K@�GbQ  �       �                   �7@@�0�!��?"            �I@ GbQ  �       �                    �?      �?             @�GbQ  ������������������������       �                      @ 146.520������������������������       �                      @.75,,Q
1�       �                    �?��0{9�?            �G@ 9,8.404�       �                    �?�X�<ݺ?             2@,0,0,37�       �                 �|Y?@��S�ۿ?             .@GbQ  �       �                 �|Y;@�����H�?             "@ 5bQ  ������������������������       �                     �?5bQ  �       �                 ���@      �?              @ 88bQ  ������������������������       �                     @ ,male,4�       �                 p&�@      �?             @8GbQ  ������������������������       ��q�q�?             @�FbQ  ������������������������       �                     �?�FbQ  ������������������������       �                     @GbQ  ������������������������       �                     @ [3bQ  �       �                  ��@V�a�� �?             =@ \GbQ  ������������������������       �                     @ ,24,0,0�       �                    �?���!pc�?             6@�FbQ  �       �                 X��A@����X�?             5@hn Henr�       �                   @'@ҳ�wY;�?	             1@�GbQ  ������������������������       �      �?             0@lip",ma������������������������       �                     �?female,������������������������       �                     @a",fema������������������������       �                     �?@�GbQ  ������������������������       �                     @ s. Albi�       �                   �0@��O���?q            @e@  GbQ  �       �                 pf�@      �?             @  Victor������������������������       �                     �? acken, �       �                    �?���Q��?             @ George�       �                 pFD!@      �?             @ �GbQ  ������������������������       �                      @Maxfiel������������������������       �                      @ Ivar S������������������������       �                     �?0IGbQ  �                         @@@���C"��?l            �d@[GbQ  �                          �? �	.��?V            ``@ahlstro�                       �!&B@�|K��2�?U             `@bre, Mi�                       �|�=@�[|x��?S            �_@�GbQ  �                       �|Y=@@-�_ .�?K            �[@75,C83,�                          �?�F��O�?7            @R@.775,,S�       �                   �:@�U�=���?1            �P@GbQ  �       �                 @3�@@9G��?'            �H@077,31.������������������������       �                     :@�,GbQ  �       �                 0S5 @���}<S�?             7@ �FbQ  �       �                   �2@      �?              @ ,44,1,0������������������������       �                     �?,female�       �                   �3@؇���X�?             @ �GbQ  ������������������������       ��q�q�?             @ Henry",������������������������       �                     @ �FbQ  ������������������������       �                     .@erine ""                       pf� @@�0�!��?
             1@. Regin������������������������       �                     "@                             ���)@      �?              @                               �;@      �?             @        ������������������������       �                      @                                �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        	                         5@؇���X�?             @        
                      �Y�@      �?              @        ������������������������       �                     �?� ��q� ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@                                �?@������?             .@                                �>@      �?              @                              (Se!@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                              pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?؇���X�?             @                             ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �        	             1@        �t�b�(z      h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �d@     �f@     �P@     �Z@     �D@     �Y@      @              A@     �Y@              3@      A@      U@      3@      ?@      *@      ,@               @      *@      @      "@      @       @              @      @      @              @      @              @      @      �?       @               @      �?       @                      �?      @              @      1@       @      .@              (@       @      @               @       @      �?      �?      �?              �?      �?              �?              @       @      @                       @      .@     �J@      (@      6@      "@      6@       @      &@              @       @       @              �?       @      @              @       @      @       @       @               @      @      &@       @      @       @                      @      @      @       @       @       @      �?       @                      �?              �?      @      @      �?               @      @      �?      �?              �?      �?              �?       @               @      �?              @              @      ?@              0@      @      .@               @      @      @      �?      @      �?      @              @      �?                      @       @              :@      @      6@              @      @               @      @      �?       @               @      �?              �?       @              Y@     �R@      �?      2@              ,@      �?      @              @      �?             �X@     �L@     @W@     �L@      @     �J@      @      D@              @      @      B@      @      <@       @      4@      �?       @      �?                       @      �?      2@              @      �?      &@      �?       @              @      �?       @      �?                       @              @      @       @      �?       @      �?      @      �?                      @              @       @                       @              *@      V@      @      A@              K@      @      ?@      @      @              <@      @      @      @      @                      @      6@      �?      &@              &@      �?       @              "@      �?       @      �?      @              7@              @             @q@     �U@      "@      1@              &@      "@      @      @               @      @               @       @      @       @                      @     �p@     �Q@      K@      E@     �B@      E@      @      5@      �?      3@      �?      @              @      �?                      0@      @       @      @      �?       @               @      �?              �?       @                      �?      @@      5@      @@      1@      3@      1@      "@      *@      �?      @      �?      �?      �?                      �?              @       @      @       @      @       @      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @                       @               @      $@      @      $@      @      @      @      @              �?      @      �?                      @      @                      �?      *@                      @      1@             �j@      <@     �h@      <@      E@      (@      E@      "@       @       @               @       @              D@      @      1@      �?      ,@      �?       @      �?      �?              @      �?      @              @      �?       @      �?      �?              @              @              7@      @      @              0@      @      .@      @      &@      @      $@      @      �?              @              �?                      @     @c@      0@      @      @      �?               @      @       @       @               @       @                      �?     �b@      *@     �]@      *@      ]@      *@      ]@      $@     @Z@      @     �P@      @     �N@      @     �G@       @      :@              5@       @      @       @              �?      @      �?       @      �?      @              .@              ,@      @      "@              @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?      �?      �?      �?                      �?      @              C@              &@      @      @      @      @       @      @                       @       @      �?       @                      �?      @      �?      @      �?      @      �?       @              �?                      @       @             �@@              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�BHzhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMIhuh*h-K ��h/��R�(KMI��h|�B@R         N                    �?�t����?�           8�@ in vers                           �?�9��L~�?^            �b@      U@                        `�@1@�C��2(�?)            �P@                                   �?�E��ӭ�?             2@                                  �?�8��8��?             (@     &@������������������������       �                     @      4@                        P��+@z�G�z�?             @        ������������������������       �                      @      &@	       
                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�q�q�?             @                               �&�)@���Q��?             @        ������������������������       �                     �?                                  �-@      �?             @        ������������������������       �                      @                                ���,@      �?              @        ������������������������       �                     �?      .@������������������������       �                     �?      @������������������������       �                     �?                                  �H@@��8��?             H@      @������������������������       �                     D@      �?                           �?      �?              @      ,@                           �?      �?             @    �L@                        ,w�U@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                     @       @       -                 pF�#@�t����?5            @U@      @       "                   �5@�#-���?            �A@      *@        !                 �{@      �?              @      @������������������������       �                     �?        ������������������������       �                     �?       @#       $                 ���@�FVQ&�?            �@@        ������������������������       �                     ,@      @%       (                 �|Y=@�KM�]�?             3@      �?&       '                   @@      �?             @     @������������������������       �                     @       ������������������������       �                     �?      @)       ,                   @@��S�ۿ?
             .@      �?*       +                 �|�=@z�G�z�?             @       ������������������������       �      �?             @      @������������������������       �                     �?       @������������������������       �                     $@      �?.       I                     @� �	��?             I@       /       D                     �?�D����?             E@     �?0       C                   �H@X�<ݚ�?             B@       1       2                 �|Y<@���!pc�?             6@       @������������������������       �                     @        3       >                    �?ҳ�wY;�?             1@     @4       ;                 `f�A@�q�q�?             (@       5       :                 X�,@@      �?              @     �?6       7                 �ܵ<@���Q��?             @        ������������������������       �                     �?      @8       9                 ��2>@      �?             @      �?������������������������       �                     @        ������������������������       �                     �?      @������������������������       �                     @      �?<       =                 @�Cq@      �?             @       ������������������������       �                     @      "@������������������������       �                     �?        ?       @                   @H@z�G�z�?             @       @������������������������       �                     �?      �?A       B                    �?      �?             @       @������������������������       �                     @        ������������������������       �                     �?      �?������������������������       �                     ,@      @E       F                 ���@@r�q��?             @     �?������������������������       �                     @      �?G       H                    �?      �?              @      @������������������������       �                     �?        ������������������������       �                     �?        J       M                    �?      �?              @        K       L                   �3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       �                   �3@�钹H��?^           ��@        P       �                    @��o	��?D             ]@       Q       v                    �?8�$�>�?4            �U@       R       S                    �?
;&����?             G@        ������������������������       �                     @        T       q                    6@�G��l��?             E@       U       n                    �?���Q��?            �A@       V       ]                    �?J�8���?             =@        W       X                   �1@z�G�z�?             @        ������������������������       �                     �?        Y       \                 ��!@      �?             @       Z       [                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ^       a                     @      �?             8@        _       `                   �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        b       g                   �1@���y4F�?             3@        c       f                   �0@      �?              @        d       e                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        h       m                 0S5 @���!pc�?             &@        i       j                   �2@      �?             @        ������������������������       �                      @        k       l                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       p                   �2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        r       s                     �?؇���X�?             @        ������������������������       �                     �?        t       u                   �1@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        w       ~                    �?z�G�z�?             D@        x       y                     @�t����?             1@       ������������������������       �                     $@        z       {                    �?����X�?             @        ������������������������       �                     @        |       }                 `f7@      �?             @       ������������������������       �                      @        ������������������������       �                      @               �                    )@��+7��?             7@       �       �                    �?�KM�]�?             3@       ������������������������       �                     *@       �       �                    �?�q�q�?             @i6bQ  �       �                    �?z�G�z�?             @ w6bQ  ������������������������       �                     @76bQ  �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @ a6bQ  �       �                    �?z�G�z�?             >@ 26bQ  �       �                    @ҳ�wY;�?             1@        ������������������������       �                     @@;6bQ  �       �                    *@��
ц��?             *@       �       �                    @�z�G��?             $@        �       �                    @      �?             @        ������������������������       �                     �?       ������������������������       �                     @t6bQ  ������������������������       �                     @        ������������������������       �                     @       ������������������������       �        	             *@        �       �                     @�/e�U��?           �{@ 6bQ  �       �                    �?      �?v             g@�6bQ  �       �                    �?*��w\��?\            �b@        �       �                    :@=QcG��?            �G@ L6bQ  �       �                   �3@���Q��?             @        ������������������������       �                      @�<6bQ  ������������������������       �                     @        �       �                   �B@�Ń��̧?             E@�3bQ  ������������������������       �                     9@       �       �                   @C@�IєX�?             1@        ������������������������       �                     �? �6bQ  ������������������������       �        
             0@        �       �                    �?��[�8��?B            �Y@        ������������������������       �                     �? �4bQ  �       �                     �?�C+����?A            @Y@       �       �                    �?���Q �?!            �H@       �       �                   �B@�z�G��?             D@       �       �                   �A@���Q��?             >@�3bQ  �       �                   �>@�q�q�?             ;@       �       �                   @>@և���X�?             5@       �       �                 �̌*@�q�q�?             2@        ������������������������       �                     @ �6bQ  �       �                 `fF<@և���X�?
             ,@       �       �                   @L@�eP*L��?             &@�4bQ  �       �                    H@      �?              @       �       �                 �|�<@      �?             @ U6bQ  ������������������������       �                     �? �6bQ  �       �                 �|�?@���Q��?             @        ������������������������       �                     �?        �       �                   �C@      �?             @ 6bQ  ������������������������       �                     �? �6bQ  ������������������������       ��q�q�?             @ �4bQ  ������������������������       �                      @        ������������������������       �                     @n6bQ  �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @��6bQ  ������������������������       �                     �?        ������������������������       �                     @ �3bQ  ������������������������       �                     @ �3bQ  ������������������������       �                     @        ������������������������       �                     $@ U6bQ  �       �                    =@X�<ݚ�?             "@ e6bQ  ������������������������       �                     �?6bQ  �       �                 ��<R@      �?              @�4bQ  �       �                   �C@z�G�z�?             @        ������������������������       �                      @        �       �                  x#J@�q�q�?             @ =/bQ  ������������������������       �                     �?6bQ  �       �                 �K@      �?              @        ������������������������       �                     �?       ������������������������       �                     �? S1bQ  ������������������������       �                     @��6bQ  �       �                    ,@4��?�?              J@d6bQ  �       �                 `f�)@�חF�P�?             ?@        ������������������������       �        	             (@ 16bQ  �       �                   �A@�d�����?             3@        �       �                 �|Y<@      �?              @ z6bQ  ������������������������       �                      @ 86bQ  �       �                 �|�=@�q�q�?             @ }6bQ  ������������������������       �                     �?       �       �                    @@���Q��?             @        ������������������������       �                     �?       ������������������������       �      �?             @       �       �                   �F@�C��2(�?             &@,6bQ  �       �                   @D@z�G�z�?             @ 5bQ  ������������������������       �                      @05bQ  ������������������������       ��q�q�?             @ �3bQ  ������������������������       �                     @        ������������������������       �                     5@``6bQ  �       �                   �M@��R[s�?            �A@�4bQ  �       �                    F@     ��?             @@6bQ  �       �                    B@�+e�X�?             9@+6bQ  �       �                    �?R���Q�?             4@W3bQ  ������������������������       �                     1@0�3bQ  ������������������������       �                     @        �       �                    �?���Q��?             @ &6bQ  ������������������������       �                      @        ������������������������       �                     @ �6bQ  ������������������������       �                     @       ������������������������       �                     @       �                          �?�����D�?�            @p@        �                          �?�ʻ����?.             Q@z6bQ  �       �                 ��@�~8�e�?$            �I@        �       �                    �?@�0�!��?             1@'6bQ  �       �                 ���@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 pff@����X�?             @|6bQ  �       �                 �|�9@      �?             @        ������������������������       �                      @        ������������������������       �                      @ �3bQ  ������������������������       �                     @ �3bQ  �       �                    �?�ʻ����?             A@        ������������������������       �                     @       �                         �>@d��0u��?             >@7bQ  �       �                 ��&@l��
I��?             ;@       �       �                   �@�r����?
             .@        �       �                 �&B@      �?             @C6bQ  �       �                   �7@�q�q�?             @        ������������������������       �                     �?T6bQ  ������������������������       �                      @ !6bQ  ������������������������       �                     �?        ������������������������       �                     &@        �                          4@      �?             (@�6bQ  �       �                   �:@      �?              @        ������������������������       �                     �?6bQ  �                           �?؇���X�?             @        ������������������������       �                     @                                �.@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              �|�:@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        	      D                ���5@     ��?v             h@       
      ?                   �?�L���?r             g@             6                ���"@d#,����?e            �d@z  �q�                          �?@�+9\J�?Z            �b@                              �|Y=@؇���X�?             5@                               ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              X�I@�KM�]�?             3@                             ���@�t����?             1@        ������������������������       �                      @                              ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @                                �7@����?K            @`@        ������������������������       �                    �A@                              ���@<����?7            �W@        ������������������������       �        	             2@                                @8@�s�c���?.            @S@                              03@      �?             @        ������������������������       �                      @        ������������������������       �                      @               1                @3�@�F��O�?,            @R@       !      "                �|Y=@X�EQ]N�?            �E@        ������������������������       �                     .@        #      0                  �C@�>4և��?             <@       $      %                pf�@�E��ӭ�?             2@        ������������������������       �                     @        &      /                   B@�q�q�?
             (@       '      .                  @@@���|���?	             &@       (      )                  �@���Q��?             $@        ������������������������       �                     @        *      +                �|�>@؇���X�?             @        ������������������������       �                     @        ,      -                �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        2      5                �|Y<@(;L]n�?             >@        3      4                  �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        7      <                �|�=@d}h���?             ,@       8      9                  �<@�C��2(�?	             &@       ������������������������       �                     @        :      ;                �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =      >                  �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @      C                pf� @P���Q�?             4@        A      B                ��Y@      �?              @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �        	             (@       E      H                   �?և���X�?             @        F      G                   �?���Q��?             @        ������������������������       �                      @       ������������������������       �                     @       ������������������������       �                      @       �t�bh�h*h-K ��h/��R�(KMIKK��h]�B�       �z@     �q@     �P@     @U@      @      N@      @      *@      �?      &@              @      �?      @               @      �?       @      �?                       @      @       @      @       @              �?      @      �?       @              �?      �?              �?      �?              �?              �?     �G@              D@      �?      @      �?      @      �?       @      �?                       @              �?              @      N@      9@      @@      @      �?      �?      �?                      �?      ?@       @      ,@              1@       @      @      �?      @                      �?      ,@      �?      @      �?      @      �?      �?              $@              <@      6@      9@      1@      4@      0@      @      0@              @      @      &@      @      @       @      @       @      @      �?              �?      @              @      �?                      @      @      �?      @                      �?      �?      @              �?      �?      @              @      �?              ,@              @      �?      @              �?      �?              �?      �?              @      @      @       @               @      @                      @     `v@     @i@      K@      O@      >@      L@      6@      8@              @      6@      4@      5@      ,@      3@      $@      �?      @              �?      �?      @      �?      �?              �?      �?                       @      2@      @      @       @      @                       @      .@      @      @      �?       @      �?      �?              �?      �?      @               @      @      �?      @               @      �?      �?      �?                      �?      @               @      @       @                      @      �?      @              �?      �?      @      �?                      @       @      @@       @      .@              $@       @      @              @       @       @               @       @              @      1@       @      1@              *@       @      @      �?      @              @      �?      �?      �?                      �?      �?              @              8@      @      &@      @      @              @      @      @      @      �?      @      �?                      @      @                      @      *@              s@     �a@      W@      W@     �T@     �P@      @      F@       @      @       @                      @      �?     �D@              9@      �?      0@      �?                      0@      T@      6@      �?             �S@      6@      @@      1@      <@      (@      2@      (@      2@      "@      (@      "@      (@      @      @               @      @      @      @      @      @      @      @              �?      @       @      �?               @       @              �?       @      �?               @      @               @      �?       @                      �?              @      @                      @      $@              @      @              �?      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                      @     �G@      @      :@      @      (@              ,@      @      @      @       @               @      @              �?       @      @      �?              �?      @      $@      �?      @      �?       @               @      �?      @              5@              "@      :@      @      :@      @      3@      @      1@              1@      @              @       @               @      @                      @      @             �j@      H@      C@      >@      6@      =@      @      ,@      �?      "@      �?                      "@       @      @       @       @               @       @                      @      3@      .@              @      3@      &@      3@       @      *@       @       @       @       @      �?              �?       @                      �?      &@              @      @       @      @      �?              �?      @              @      �?      @      �?                      @      @                      @      0@      �?              �?      0@             �e@      2@     @e@      .@     �b@      ,@     �a@      &@      2@      @      �?      �?      �?                      �?      1@       @      .@       @       @              @       @      @       @      �?               @             �^@       @     �A@             �U@       @      2@             @Q@       @       @       @               @       @             �P@      @      C@      @      .@              7@      @      *@      @      @              @      @      @      @      @      @              @      @      �?      @               @      �?      �?              �?      �?      �?                      �?      $@              =@      �?       @      �?       @                      �?      ;@              &@      @      $@      �?      @              @      �?              �?      @              �?       @               @      �?              3@      �?      @      �?      @                      �?      (@              @      @       @      @       @                      @       @        �t�bubhhubehhub.